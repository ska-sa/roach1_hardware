* AD711T SPICE Macro-model       		1/91, Rev. A
*								JLW / PMI
*
* This version of the AD711 model simulates the worst case
* parameters of the 'T' grade. The worst case parameters 
* used correspond to those in the data book.
*
*
* Copyright 1991 by Analog Devices, Inc.
*
* Refer to "README.DOC" file for License Statement.  Use of this model
* indicates your acceptance with the terms and provisions in the License Statement.
*
* connections:  non-inverting input 
*               |  inverting input  
*               |  |  positive supply
*               |  |  |  negative supply
*               |  |  |  |  output
*               |  |  |  |  |
.SUBCKT AD711T 13 15 12 16 14
* 
VOS 15 8 DC 0.5E-3
EC 9 0 (14,0) 1
C1 6 7 .5E-12
RP 16 12 10.35E3
GB 11 0 (3,0) 1.67E3
RD1 6 16 16E3
RD2 7 16 16E3
ISS 12 1 DC 100E-6
CCI 3 11 45E-12
GCM 0 3 (0,1) 1.76E-9
GA 3 0 (7,6) 780E-6
RE 1 0 2.5E6
RGM 3 0 2.6E3
VC 12 2 DC 2.8
VE 10 16 DC 3.1
RO1 11 14 25
CE 1 0 2E-12
RO2 0 11 30
RS1 1 4 5.77E3
RS2 1 5 5.77E3
J1 6 13 4 FET
J2 7 8 5 FET
DC 14 2 DIODE
DE 10 14 DIODE
DP 16 12 DIODE
D1 9 11 DIODE
D2 11 9 DIODE
IOS 15 13 12.5E-12
.MODEL DIODE D()
.MODEL FET PJF(VTO=-1 BETA=1E-3 IS=50E-12)
.ENDS
