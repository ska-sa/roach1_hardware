* OP221E SPICE Macro-model                 9/91, Rev. A
*                                           JCB / PMI
*
* This version of the OP-221 model simulates the worst case 
* parameters of the 'E' grade.  The worst case parameters
* used correspond to those in the data sheet.
*
* Copyright 1991 by Analog Devices, Inc.
*
* Refer to "README.DOC" file for License Statement.  Use of this model
* indicates your acceptance with the terms and provisions in the License Statement.
*
* Node assignments
*                non-inverting input
*                | inverting input
*                | | positive supply
*                | | |  negative supply
*                | | |  |  output
*                | | |  |  |
.SUBCKT OP221E   1 2 99 50 31
*
* INPUT STAGE & POLE AT 1.9 MEGHZ
*
R1    2  3     5E11
R2    1  3     5E11
R3    5 50     5160
R4    6 50     5160
CIN   1  2     2E-12
C2    5  6     8.12E-12
I1    99 4     10E-6
IOS   1  2     1.5E-9
EOS   9  1     POLY(1)  24 27  150E-6  1
Q1    5  2  4  QX
Q2    6  9  4  QX
*
EREF  98 0     27  0  1
*
* FIRST GAIN STAGE
*
R5   10 98     1E6
G1   98 10     5  6  39E-6
D1   10 11     DX
D2   12 10     DX
E1   99 11     POLY(1) 99 27 -1.4 1
E2   12 50     POLY(1) 27 50 -1.4 1
*
* GAIN STAGE & DOMINANT POLE AT 0.41 HZ
*
R7   13 98     7.7E9
C3   13 98     50E-12
G2   98 13     10  27  5E-6
V1   99 14     1.45
V2   15 50     1.3
D3   13 14     DX
D4   15 13     DX
*
* POLE AT 3.0 MEGHZ
*
R8   16 98     1E6
C5   16 98     53.1E-15
G3   98 16     13 27  1E-6
*
* POLE AT 3.0 MEGHZ
*
R9   17 98     1E6
C7   17 98     53.1E-15
G10  98 17     16 27  1E-6
*
* COMMON-MODE GAIN NETWORK WITH ZERO AT 31.6 HZ
*
R10  24 98     1
R11  23 24     1E6
C4   23 24     5.033E-9
E4   98 23     3  27  31.62
*
* POLE AT 3.0 MEGHZ
*
R12  25 98     1E6
C6   25 98     53.1E-15
G9   98 25     17 27  1E-6
*
* OUTPUT STAGE
*
ISY  99 50     290E-6
R13  27 99     150E3
R14  27 50     150E3
R15  30 99     450
R16  30 50     450
L1   30 31     1E-8
G4   28 50     25 30  2.22E-3
G5   29 50     30 25  2.22E-3
G6   30 99     99 25  2.22E-3
G7   50 30     25 50  2.22E-3
D5   99 28     DX
D6   99 29     DX
D7   50 28     DY
D8   50 29     DY
D9   25 33     DX
V3   33 30     1.6
D10  32 25     DX
V4   30 32     1.6
*
* MODELS USED
*
.MODEL QX PNP(BF=63.7)
.MODEL DX   D(IS=1E-15)
.MODEL DY   D(IS=1E-15 BV=50)
.ENDS
