* ADN8830 Long-Time SPICE Model v0.3
* 
* Copyright 2001 Analog Devices, Inc.
* TAM 12/01
*
* Note: This model is for long time (>100ms) transient reponse simulations
*       of the entire ADN8830-TEC-Object-Thermistor loop.  To speed up
*       simulation it does not use external transistors, instead driving the
*       TEC directly from Pins 9 and 19.
*
* Note: Node numbers 1-32 refer to actual pin numbers on device
*
*		  THERMFAULT
*		  | THERMIN
*		  | | TEMPSET
*		  | | | TEMPLOCK
*		  | | | | 1.5V
*		  | | | | | VREF
*		  | | | | | | AVDD
*		  | | | | | | | OUT_B
*		  | | | | | | | |  TEMPCTL
*		  | | | | | | | |  |  COMPFB
*		  | | | | | | | |  |  |  COMPOUT
*		  | | | | | | | |  |  |  |  OUT_A
*		  | | | | | | | |  |  |  |  |  PVDD
*		  | | | | | | | |  |  |  |  |  |  PGND
*		  | | | | | | | |  |  |  |  |  |  |  AGND
*		  | | | | | | | |  |  |  |  |  |  |  |  TEMPOUT
*		  | | | | | | | |  |  |  |  |  |  |  |  |
.SUBCKT ADN8830_L 1 2 4 5 6 7 8 9 12 13 14 19 20 23 30 31
*
* Reference voltages
*
V15  6 30 1.5V
V30 33 30 3.0V
*
* THERMFAULT Output
*
V6 71 30 2.3V
V7 72 30 0.2V
O4  2 71 ADCONV  DGTLNET=54  IO_CMOS
O5 72  2 ADCONV  DGTLNET=55  IO_CMOS
U8 OR(2) 8 30 54 55 56 T_STD IO_CMOS
N5  1 30 8 DACONV DGTLNET=56 IO_CMOS
*
* TEMPLOCK Output
*
V8 73 30 1.55V
V9 74 30 1.45V
O6 73 12 ADCONV DGTLNET=57    IO_CMOS
O7 12 74 ADCONV DGTLNET=58    IO_CMOS
U9 AND(2) 8 30 57 58 59 T_STD IO_CMOS
N6  5 30  8 DACONV DGTLNET=59 IO_CMOS
*
* Output Amplifiers
*
EOUTB  96  6 (14,6) -14
EOUTA  97 23 POLY(2) (14,6) (9,23) 0 4 1

ELIN  9 23 VALUE={LIMIT( V(96), V(23), V(20) )}
EPWM 19 23 VALUE={LIMIT( V(97), V(23), V(20) )}

*
* Compensation Amplifier
*
* E1    95 30 (6,93) 100k
* RD1   95 30 1
* ECOMP 98 30 VALUE={LIMIT( V(95), V(30), V(33) )}
* RD2   98 30 1
* RD3   12 93 100k
* RD4   93 98 100k

X2  6 13 14 33 30 OPAMP
*
* Input Error Amplifier
*
E2 34  6 POLY(1) (4,2) 0 20 ; (TEMPSET-THERMIN)*20 + 1.5V
X3 34 12 12 33 30 OPAMP

VREF 7 30 2.45V
*
* TEMPOUT Amplifier
*
E3  35  6 (4,2) 3
R10 35 31 0.1
*
.MODEL ADCONV DOUTPUT(RLOAD=1E8,S0NAME="0",S0VLO=-10,S0VHI=0,
+                               S1NAME="1",S1VLO=0,S1VHI=10)
.MODEL T_STD UGATE()
.MODEL DACONV DINPUT(S0NAME="0",S0TSW=20ns,S0RLO=2,S0RHI=5E6,
+                    S1NAME="1",S1TSW=20ns,S1RLO=5E6,S1RHI=2,
+                    S2NAME="X",S2TSW=20ns,S2RLO=5E6,S2RHI=5E6,
+                    S3NAME="Z",S3TSW= 1ns,S3RLO=5E6,S3RHI=5E6)
.MODEL IO_CMOS UIO()
.MODEL DX D(IS=1E-14,RS=1m)
.ENDS
*
* Simple Op Amp Avo=120k
*
.SUBCKT OPAMP 1 2 3 99 50
G1 50  4 (2,1) 1
R1  4 50 100k
C1  4 50 1.5p
D1  4 98 DX
V1 99 98 0.6
D2 51  4 DX
V2 51 50 0.6
M1  3  4 50 50 NAMPFET L=1u W=10m
R2 99  3 10k
.MODEL DX D(IS=1E-14,RS=1m)
.MODEL NAMPFET NMOS(LEVEL=1,VTO=0,KP=24E-6)
.ENDS
*$