*	AD8062 SPICE 
*				MACRO MODEL REV 0
*						M.M 9/4/02
*This model will give the typical performance characteristics
*for the following parameters:

*************************************************************
*	Bandwidth
*	Slewrate
*	Open Loop Gain/Phase
*	Supply Currents
*	Output current should reflect back to the supplies
*	Output current (short circuit limiting)
*	Output resistance (dc)
*	Input voltage range
*	Output voltage range
*  Vos is static and will not vary
*  CMRR is not modeled
*  Distortion is not characterized
************************************************************

* Node assignments |Non-Inverting input	
*		   |	|Inverting input			
*		   |	|	|Positive supply
*		   |	|	|	|Negative supply
*		   |	|	|	|	|Output
*		   |	|	|	|	|
.SUBCKT AD8062 	   1	2	99	50      45
* Input stage *

I1 4 50 1.25E-3
Q1 5 2 10 QPI 	
Q2 6 9 11 QPI
Vos 9 1 0
*IOS 2 1 .3u
R1 1 3 6.5e6
R2 3 2 6.5e6
Cin 2 1 1p
R3 99 5 2.5k
R4 99 6 2.5k
R5 10 4 948
R6 11 4 948
*C  5 6 .16p


*Gain and Pole stage w/ pole at 17 kHz*

Eref 98 0 POLY(2) 99 0 50 0 0 .5 .5 

R7  12 98 6.04e6
C2  12 98 1.54pf
G1  98 12 5 6 6.54e-4
v1 99 14 -.95
v2 16 50 -.95
D1 12 14 Dx
D2 16 12 Dx

*Zero at 90 MHz and pole at 500*
Gzp  98 25 12 98 .92
Rzp2 25 26 6.5
Rzp1 26 98 1
Lzp 25 26 1.72e-9


*pole at 500 MHz
G2 98 27 25 98 .85
Rp3 98 27 1
Cp 98 27 318p


*Eout 32 98 25 98 1
*Rout 33 32 .17



*Buffer Stage
Gbuf 98 32 27 98 1e-2
Rbug 32 98 100

* COMMON-MODE GAIN NETW0RK
Ecm 20 98 POLY(2) 2 98 1 98 0 .5 .5 
Gcm 98 21 20 98 .4e-6
L4 21 23 1e-3
Rx 23 98 1k


*Output Stage *
R8 99 33 .17
R9 33 50 .17
G23 33 99 99 32 5.88
G24 50 33 32 50 5.88
G25 98 52 33 32 5.88
D7 52 53 Dx
D8 54 52 Dx
V8 53 98 0
V9 98 54 0
V6  34 33 -.849
V7  33 35 -.849
D5  32 34 Dx
D6  35 32 Dx
Vcd 45 33 0


Fol 98 72 vcd 1
Vi1 72 70 0
Vi2 72 71 0
D11 70 98 Dx
D12 98 71 Dx

Erefq 96 0 45 0 1
Fq1 99 96 POLY(2) Vi2 Vcd 0 1 -1
Fq2 96 50 POLY(2) Vi1 Vcd 0 1 -1



* Quiescent Current

Ibias 99 50 -5.15m


.MODEL d1 D(IS=10e-15)
.MODEL Dy D(IS=10e-15)
.MODEL Dx D(IS=10e-15)
.MODEL Dz D(IS=10e-15)
.MODEL QPI NPN(IS=100e-18 NF=1 BF=178.4)
.ENDS








