* AD8067 Spice Model  Rev. A, 3/2004 TRW
*
* Refer to "README.DOC" file for License Statement.
* Use of this model indicates your acceptance with
* the terms and provisions in the License Statement.
*
* The following parameters are accurately modeled;
*
*       Open loop gain and phase vs. frequency
*       Output impedance vs. frequency
*       Output clamping voltage and current
*       FET Input common mode range
*       Voltage noise
*       Output currents are reflected to V supplies
*       Vos is static and will not vary
*       Distortion is not characterized       
*
*
*    Node assignments
*              non-inverting input
*              | inverting input
*              | | positive supply
*              | | |  negative supply
*              | | |  |  output
*              | | |  |  |
.SUBCKT AD8067 1 2 99 50 45

* FET INPUT STAGE

Eos 9 2 poly(1) 100 98 39m 1
Cd 1 2 2.5p
Ccm1 1 0 1.5p
Ccm2 2 0 1.5p
J1 5 1 4 pmod 
J2 6 9 4 pmod
Ib1 1 0 5.6p
Ib2 9 0 5.6p
R3 50 5 rnoise 1
R4 50 6 rnoise 1
I11 99 4 1
*R5 73 4 390
*R6 74 4 390

* Common Mode Clamp

Vcmc 99 77 5.65
Dcmc 4 77 dx

* COMMON-MODE GAIN NETW0RK

Ecm 80 98 POLY(2) 2 98 1 98 0 .5 .5 

* GAIN STAGE & POLE AT 400Hz

Ecc 97 0 99 0 1
Ess 52 0 50 0 1
Eref 98 0 POLY(2) 99 0 50 0 0 .5 .5 

G1 13 98 5 6 .0035e3
R7 13 98 Rnoise 255e3
C3 13 98 1.56e-9
V1 97 14 0.7
V2 16 52 0.75
D1 13 14 DX
D2 16 13 DX

* POLE AT 60 MHz
G2 98 43 13 98 1
R10 98 43 rnoise 1
C5 98 43 2.65n

* POLE AT 130 MHz
G3 98 53 43 98 1
R11 98 53 rnoise 1
C6 98 53 1.22n

*POLE AT 130 MHz
G4 98 63 53 98 1
R12 98 63 rnoise 1
C7 98 63 1.22n

* BUFFER STAGE
Gbuf 98 81 63 98 1e-2
Rbuf 81 98 Rnoise 100
* OUTPUT STAGE

Vo1 99 90 0
Vo2 51 50 0
R18 25 90 rnoise .02
R19 25 51 rnoise .02
Vcd 25 45 0
G6 25 90 99 81 50
G7 51 25 81 50 50
V4 26 25 -0.838
V5 25 27 -0.838
D5 81 26 Dx
D6 27 81 DX

Fo1 98 70 vcd 1
D7 70 71 DX
D8 72 70 DX
vi1 71 98 0
Vi2 98 72 0

Erefq 96 0 45 0 1 
Iq 99 50 -0.1017
Fq1 96 99 POLY(2) Vo1 Vi1 0 1 -1
Fq2 50 96 POLY(2) Vo2 Vi2 0 1 -1

****** Voltage noise stage

rnoise1 39 98 5.5e-4
vnoise1 39 98 0
vnoise2 101 98 0.75
dnoise1 101 39 dn
fnoise1 100 98 vnoise1 1
rnoise2 100 98 1

.model Rnoise RES(T_abs=-373)
.model pmod pjf beta=1e-2
.MODEL DX D
.model dn d(kf=2e-12,af=1)

.ENDS
