* AD680 SPICE Macromodel 5/94, Rev. A
* AAG / ADSC
*
* Copyright 1994 by Analog Devices, Inc.
*
* Refer to "README.DOC" file for License Statement.  
* Use of this model indicates your acceptance with 
* the terms and provisions in the License Statement.
*
*  NODE NUMBERS
*              VIN
*              |  TEMP
*              |  |  GND
*              |  |  |  VOUT
*              |  |  |  |
.SUBCKT AD680  2  3  4  6
*
* BANDGAP REFERENCE
*
IBG 4 10 DC 1.2864651E-3
RBG 10 4 1E3 TC=10E-6
EN 10 11 14 0 1
G1 4 11 2 4 2.0584285E-8
F1 4 11 VLR 4.116857E-5
Q1 2 11 12 QT
I1 12 4 DC 50E-6
R1 12 3 11.486E3
I2 3 4 DC 0
*
* NOISE VOLTAGE GENERATOR
*
VN1 13 0 DC 2
DN1 13 14 DEN
DN2 14 15 DEN
VN2 0 15 DC 2
*
* INTERNAL OP AMP AND DOMINANT POLE @ 0.2 Hz
*
G2 4 16 11 24 2.513274E-4
R2 16 4 7.957747E9
C1 16 4 1E-10
D1 16 17 DX
V1 2 17 DC 1.3
*
* SECONDARY POLE @ 300 kHz
*
G3 4 18 16 4 1E-6
R3 18 4 1E6
C2 18 4 5.3051647E-13
*
* OUTPUT STAGE
*
ISY 2 4 8.693E-5
FSY 2 4 V1 -1
RSY 2 4 2.5E6
*
G4 4 21 18 4 1E-3
R4 21 4 1E3
FSC 21 4 VSC 1
VSC 2 19 DC 0
Q2 19 2 20 QN
RSC 2 20 26
Q3 20 21 22 QN
R5 22 24 21.6E3
R6 24 4 22.9E3
VLR 23 22 DC 0
L1 23 6 1E-7
*
.MODEL QT NPN(IS=1.5E-16 BF=1E3 XTI=7.2)
.MODEL QN NPN(IS=1E-15 BF=1E3)
.MODEL DX D(IS=1E-15)
.MODEL DEN D(IS=1E-12 RS=1.98709E+06 AF=1 KF=1.21245E-16)
.ENDS AD680
