***** AD8023 SPICE model       Rev A SMR/ADI 7-14-97

* Copyright 1997 by Analog Devices, Inc.

* Refer to "README.DOC" file for License Statement.  Use of this model
* indicates your acceptance with the terms and provisions in the License Statement.

* This model will give typical performance characteristics
* for the following parameters;

*     closed loop gain and phase vs bandwidth
*     output current and voltage limiting
*     offset voltage (is static, will not vary with vcm)
*     ibias (again, is static, will not vary with vcm)
*     slew rate and step response performance
*     (slew rate is based on 10-90% of step response)
*     current on output will be reflected to the supplies 
*     vnoise, referred to the input
*     inoise, referred to the input

*     distortion is not characterized

* Node assignments
*                non-inverting input
*                | inverting input
*                | | positive supply
*                | | |  negative supply
*                | | |  |  output
*                | | |  |  |
.SUBCKT AD8023an 1 2 99 50 28

* input stage *

q1 50 3 5 qp1
q2 99 5 4 qn1
q3 99 3 6 qn1
q4 50 6 4 qp1
i1 99 5 173e-6
i2 6 50 173e-6
cin1 1 98 2e-12
cin2 2 98 2e-12
v1 4 2 0

* input error sources *

eos 3 1 poly(1) 20 98 2e-3 0
fbn 2 98 poly(1) vnoise3 10e-6 0
fbp 1 98 poly(1) vnoise3 5e-6 0

* slew limiting stage *

fsl 98 16 v1 1
dsl1 98 16 d1
dsl2 16 98 d1
dsl3 16 17 d1
dsl4 17 16 d1
rsl  17 18 3.5
vsl  18 98 0

* gain stage *

f1 98 7 vsl 2
rgain 7 98 2e5
cgain 7 98 1.7e-12
dcl1 7 8 d1
dcl2 9 7 d1
vcl1 99 8 1.7
vcl2 9 50 1.7
           
* second pole *

epole1 14 98 7 98 1
rpole1 14 15 1
*cpole1 15 98 2.5e-10
cpole1 15 98 2e-10

* third pole *

epole2 34 98 15 98 1
rpole2 34 35 1
*cpole2 35 98 2.5e-10
cpole2 35 98 2e-10

* reference stage *

eref 98 0 poly(2) 99 0 50 0 0 0.5 0.5 

ecmref 30 0 poly(2) 1 0 2 0 0 0.5 0.5

* vnoise stage *

rnoise1 19 98 1.84e-3
vnoise1 19 98 0
vnoise2 21 98 0.53
dnoise1 21 19 dn

fnoise1 20 98 vnoise1 1
rnoise2 20 98 1

* inoise stage *

rnoise3 22 98 8.18e-6
vnoise3 22 98 0
vnoise4 24 98 0.575
dnoise2 24 22 dn

fnoise2 23 98 vnoise3 1
rnoise4 23 98 1

* buffer stage *

gbuf 98 13 35 98 1e-2
rbuf 98 13 1e2

* output current reflected to supplies *

fcurr 98 40 voc 1
vtest 40 25 0
vcur1 25 26 0
vcur2 27 25 0
dcur1 26 98 d1
dcur2 98 27 d1
fsy 99 50 poly(2) vcur1 vcur2 9.2e-3 0 0

* output stage *

gout1 99 10 13 99 0.5
gout2 50 10 13 50 0.5
rout1 10 99 2
rout2 10 50 2
voc 10 28 0
rout3 28 98 1e6
dcl3 13 11 d1
dcl4 12 13 d1
vcl3 11 10 -0.585
vcl4 10 12 -0.585

.model qp1 pnp()
.model qn1 npn()
.model d1  d()
.model dn  d(af=1 kf=1e-8)
.ends AD8023
