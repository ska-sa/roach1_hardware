* OP292G SPICE Macro-model              Rev. A, 3/95
*                                       ARG / ADSC
*
* This version of the OP292 model simulates the worst-case
* parameters of the 'G' grade. The worst-case parameters
* used correspond to those in the data sheet.
*
* Copyright 1995 by Analog Devices
*
* Refer to "README.DOC" file for License Statement. Use of
* this model indicates your acceptance of the terms and pro-
* visions in the License Statement.
*
* Node assignments
*                non-inverting input
*                |  inverting input
*                |  |  positive supply
*                |  |  |  negative supply
*                |  |  |  |  output
*                |  |  |  |  |
.SUBCKT OP292G   2  1  99 50 34
*
* INPUT STAGE AND POLE AT 40MHZ
*
I1   99   4    51.4E-6
IOS  2    1    25E-9
EOS  2    3    POLY(1) (21,30) 2E-3 16.8
CIN  1    2    2E-12
Q1   5    1    7    QP
Q2   6    3    8    QP
R3   5    50   2E3
R4   6    50   2E3
R5   4    7    965
R6   4    8    965
C1   5    6    .995E-12
*
* GAIN STAGE
*
EREF 98   0    (30,0) 1
G1   98   9    (5,6) 500E-6
R7   9    98   14.388E3
D1   9    10   DX
D2   11   9    DX
V1   99   10   .6
V2   11   50   .6
*
* ZERO/POLE AT 6MHZ/12MHZ
*
E1   12   98   (9,30) 2
R8   12   13   1
R9   13   98   1
C3   12   13   26.526E-9
*
* ZERO AT 15MHZ
*
E2   14   98   (13,30) 1E6
R10  14   15   1E6
R11  15   98   1
C4   14   15   10.610E-15
*
* COMMON MODE STAGE WITH ZERO AT 40KHZ
*
ECM  20   98   POLY(2) (1,30) (2,30) 0 0.5 0.5
R20  20   21   1E6
R21  21   98   10
*C5   20   21   3.979E-12
*
* POLE AT 100MHZ
*
G2   98   16   (9,30) 1
R12  16   98   1
C6   16   98   1.592E-9
*
* OUTPUT STAGE
*
RS1  99   30   1E6
RS2  30   50   1E6
ISY  99   50   .236E-3
G3   31   50   POLY(1) (16,30) -1.681511E-6 1E-6
R16  31   50   1E6
DCL  50   31   DZ
I2   99   32   250E-6
RCP  99   36   75
RCL  33   50   75
Q6   35   36   99   QPA
Q7   32   37   50   QNA
R17  35   37   1E3
M1   32   31   50   50   MN L=9E-6 W=1000E-6 AD=15E-9 AS=15E-9
M2   34   31   50   50   MN L=9E-6 W=1000E-6 AD=15E-9 AS=15E-9
CC   31   32   0.23E-12
Q3   36   32   34   QNA
Q4   33   32   34   QPA
Q5   31   33   50   QNA
.MODEL QNA NPN(IS=1.19E-16 BF=253 VAF=193 RC=400)
.MODEL QPA PNP(IS=5.21E-17 BF=131 VAF=62 RC=250)
.MODEL MN NMOS(LEVEL=3 VTO=1.3 RS=0.3 RD=0.3 LD=1.48E-6 WD=1E-6)
.MODEL QP PNP(BF=35.714)
.MODEL DX D
.MODEL DZ D(BV=3.6)
.ENDS OP292G
