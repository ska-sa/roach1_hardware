* AD633J Analog Multiplier Macro Model 12/93, Rev. A
* AAG/PMI
*
* This version of the AD633 analog multiplier model simulates the worst case
* parameters of the 'J' grade.  The worst case parameters used correspond
* to those parameters in the data sheet.
*
* Copyright 1993 by Analog Devices, Inc.
*
* Refer to "README.DOC" file for License Statement.  Use of this model
* indicates your acceptance with the terms and provisions in the License Statement.
*
* Node assignments
*              X1
*              |  X2
*              |  |  Y1
*              |  |  |  Y2
*              |  |  |  |  VNEG
*              |  |  |  |  |  Z
*              |  |  |  |  |  |  W
*              |  |  |  |  |  |  |  VPOS
*              |  |  |  |  |  |  |  |
.SUBCKT AD633J 1  2  3  4  5  6  7  8
*
EREF 100 0 POLY(2) 8 0 5 0 (0,0.5,0.5)
*
* X-INPUT STAGE & POLE AT 15 MHz
*
IBX1 1 0 DC 2E-6
IBX2 2 0 DC 2E-6
EOSX 10 1 POLY(1) (16,100) (30E-3,1)
RX1A 10 11 5E6
RX1B 11 2 5E6
*
GX 100 12 10 2 1E-6
RX 12 100 1E6
CX 12 100 1.061E-14
VX1 8 13 DC 3.05
DX1 12 13 DX
VX2 14 5 DC 3.05
DX2 14 12 DX
*
* COMMON-MODE GAIN NETWORK WITH ZERO AT 560 Hz
*
ECMX 15 100 11 100 10
RCMX1 15 16 1E6
CCMX 15 16 2.8421E-10
RCMX2 16 100 1
*
* Y-INPUT STAGE & POLE AT 15 MHz
*
IBY1 3 0 DC 2E-6
IBY2 4 0 DC 2E-6
EOSY 20 3 POLY(1) (26,100) (30E-3,1)
RY1A 20 21 5E6
RY1B 21 4 5E6
*
GY 100 22 20 4 1E-6
RY 22 100 1E6
CY 22 100 1.061E-14
VY1 8 23 DC 3.05
DY1 22 23 DX
VY2 24 5 DC 3.05
DY2 24 22 DX
*
* COMMON-MODE GAIN NETWORK WITH ZERO AT 560 Hz
*
ECMY 25 100 21 100 10
RCMY1 25 26 1E6
CCMY 25 26 2.8421E-10
RCMY2 26 100 1
*
* Z-INPUT STAGE & POLE AT 15 MHz
*
IBZ1 7 0 DC 8E-7
IBZ2 6 0 DC 8E-7
RZ1 7 6 10E6
*
GZ 100 32 7 6 1E-6
RZ2 32 100 1E6
CZ 32 100 1.061E-14
VZ1 8 33 DC 3.05
DZ1 32 33 DX
VZ2 34 5 DC 3.05
DZ2 34 33 DX
*
* 50-MHz MULTIPLIER CORE & SUMMER
*
GXY 100 40 POLY(2) (12,100) (22,100) (0,0,0,0,0.1E-6)
RXY 40 100 1E6
CXY 40 100 3.1831E-15
*
* OP AMP INPUT STAGE
*
VOOS 59 40 DC 50E-3
Q1 55 32 60 QX
Q2 56 59 61 QX
R1 8 55 3.1831E4
R2 60 54 3.1313E4
R3 8 56 3.1831E4
R4 61 54 3.1313E4
I1 54 5 1E-4
*
* GAIN STAGE & DOMINANT POLE AT 316.23 Hz
*
G1 100 62 55 56 3.141637E-5
R5 62 100 1.0066E8
C3 62 100 5E-12
V1 8 63 DC 4.3399
D1 62 63 DX
V2 64 5 DC 4.3399
D2 64 62 DX
*
* NEGATIVE ZERO AT 20 MHz
*
ENZ 65 100 62 100 1E6
RNZ1 65 66 1
FNZ 65 66 VNC -1
RNZ2 66 100 1E-6
ENC 67 0 65 66 1
CNZ 67 68 7.9577E-9
VNC 68 0 DC 0
*
* POLE AT 4 MHz
*
G2 100 69 66 100 1E-6
R6 69 100 1E6
C2 69 100 3.9789E-14
*
* OP AMP OUTPUT STAGE
*
FSY 8 5 POLY(2) VZC1 VZC2 (4.8286E-3,1,1)
RDC 8 5 28E3
GZC 100 73 72 69 11.623E-3
VZC1 74 100 DC 0
DZC1 73 74 DX
VZC2 100 75 DC 0
DZC2 75 73 DX
VSC1 70 72 1.125
DSC1 69 70 DX
VSC2 72 71 1.125
DSC2 71 69 DX
GO1 72 8 8 69 11.623E-3 
RO1 8 72 86
GO2 5 72 69 5 11.623E-3 
RO2 72 5 86
LO 72 7 1E-7
*
* MODELS USED
*
.MODEL QX NPN(BF=1E4)
.MODEL DX D(IS=1E-15)
.ENDS AD633J
