* AD745A SPICE Macro-model              10/95, Rev. B
*                                       ARG / ADSC
*
* This version of the AD745 model simulates the worst-case
* parameters of the 'A' grade. The worst-case parameters
* used correspond to those in the data sheet.
*
*
* Revision History:
*     Rev. B
* Changed the negative zero circuit to correspond to the new design
* which eliminates the negative capacitor value.
*
*
* Copyright 1992 by Analog Devices, Inc.
*
* Refer to "README.DOC" file for License Statement. Use of this model
* indicates your acceptance with the terms and provisions in the License
* Statement.
*
* Node assignments
*                non-inverting input
*                |  inverting input
*                |  |  positive supply
*                |  |  |  negative supply
*                |  |  |  |  output
*                |  |  |  |  |
.SUBCKT AD745A   3  2  99 50 37
*
* INPUT STAGE AND POLE AT 54MHZ
*
I1   97   1    1
J1   5    2    1    JX
J2   6    4    1    JX
CIN  2    3    20E-12
IOS  3    2    75E-12
EN   7    3    9 0 1
GN1  0    2    12 0 1E-6
GN2  0    3    15 0 1E-6
EOS  4    7    POLY(1) 31 52 800E-6 1
R1   5    51   86.842E-3
R2   6    51   86.842E-3
C1   5    6    16.969E-9
EPOS 97   0    99 0 1
ENEG 51   0    50 0 1
EREF 98   0    52 0 1
*
* VOLTAGE NOISE SOURCE WITH FLICKER NOISE
*
VN1  8    0    DC 2
VN2  0    10   DC 2
DN1  8    9    DEN
DN2  9    10   DEN
*
* CURRENT NOISE SOURCE WITH FLICKER NOISE
*
VN3  11   0    DC 10
VN4  0    13   DC 10
DN3  11   12   DIN
DN4  12   13   DIN
*
* CURRENT NOISE SOURCE WITH FLICKER NOISE
*
VN5  14   0    DC 10
VN6  0    16   DC 10
DN5  14   15   DIN
DN6  15   16   DIN
*
* GAIN STAGE AND DOMINANT POLE AT 22.9HZ
*
R3   17   98   86.842E3
C2   17   98   80E-9
G1   98   17   5 6 11.515
V1   97   18   .727
V2   19   51   1.893
D1   17   18   DX
D2   19   17   DX
*
* POLE AT 30MHZ
*
R4   23   98   1
C3   23   98   5.305E-9
G2   98   23   17 52 1
*
* POLE AT 30MHZ
*
R5   24   98   1
C4   24   98   5.305E-9
G3   98   24   23 52 1
*
* NEGATIVE ZERO AT -54MHZ
*
R6   25   26   1
R7   26   98   1E-6
E1   25   98   24 52 1E6
VX1  84   0    DC 0
EX1  83   0    25 26 1
FX1  25   26   VX1 -1
CX1  83   84   2.947E-9
*
* POLE / ZERO AT 2MHZ / 2.25MHZ
*
R8   27   98   1
R9   27   28   8
C6   28   98   8.842E-9
G4   98   27   26 52 1
*
* COMMON MODE GAIN STAGE WITH ZERO AT 126KHZ
*
E2   29   30   2 52 0.5
E3   30   98   3 52 0.5
R10  29   31   1
R11  31   98   100E-6
C7   29   31   1.264E-6
*
* REFERENCE NODE AND OUTPUT STAGE
*
RMP1 97   52   1
RMP2 52   51   1
GSY  99   50   POLY(1) 99 50 9.625E-3 12.5E-6
R13  99   36   200
R14  36   50   200
L1   36   37   1E-10
G5   34   50   27 36 5E-3
G6   35   50   36 27 5E-3
G7   36   99   99 27 5E-3
G8   50   36   27 50 5E-3
V3   32   36   1.55
V4   36   33   1.55
D3   27   32   DX
D4   33   27   DX
D5   99   34   DX
D6   99   35   DX
D7   50   34   DY
D8   50   35   DY
F1   36   0    V3 1
F2   0    36   V4 1
*
* MODELS USED
*
.MODEL JX PJF(BETA=66.299, VTO=-1.5 IS=400E-12)
.MODEL DX D(IS=1E-15)
.MODEL DY D(IS=1E-15, BV=50)
.MODEL DEN D(RS=1.931E3, KF=2.278E-15, AF=1)
.MODEL DIN D(RS=5.277E3, KF=42.593E-15, AF=1)
.ENDS AD745A
