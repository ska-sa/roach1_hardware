*       AD8024 Spice Model  Rev. A, 4/01
*                           VC
*
*       Copyright 2000 by Analog Devices, Inc.
*
*       Refer to "README.DOC" file for License Statement.
*       Use of this model indicates your acceptance with
*       the terms and provisions in the License Statement
*
*       The following parameters are accurately modeled
*
*       Closed loop gain and phase vs. frequency
*       Output clamping voltage and current
*       Slew rate and step response performance
*       Output currents are reflected to V supplies
*       Vos is static and will not vary
*       Input resistance adjusted to stablize amplifier
*       Distortion is not characterized       
*       Common mode rejection ratio is not modeled
*       Noise is not modeled
*
*     Node assignments
*              Non-Inverting Input
*              | Inverting Input 
*              | | positive supply
*              | | |  negative supply
*              | | |  |  output
*              | | |  |  | 
*              | | |  |  |
.SUBCKT AD8024 1 2 99 50 30
* INPUT STAGE
VL1 8 2 0
I1 99 5 3e-6
I2 4 50 3e-6
Q1 50 3 5 QP1
Q2 99 3 4 QN1
Q3 99 5 8 QN2
Q4 50 4 8 QP2

* INPUT ERROR SOURCES
IB1 99 2 1e-6
IB2 99 3 1e-6
VOS 3 1 2m
               
* SLEW RATE LIMITING STAGE
FL1 98 40 VL1 1
DL1 40 98 DX
DL2 98 40 DX
DL3 40 42 DX
DL4 42 40 DX
VL2 42 43 0
RL1 43 98 8.5k

* GAIN STAGE
Eref 98 0 POLY(2) 99 0 50 0 0 .5 .5 
F1 98 13 VL2 2
R7 98 13 1.2Meg
C3 98 13 75f
V1 99 14 2
V2 16 50 2
D1 13 14 DX
D2 16 13 DX

* 2nd POLE STAGE
G2 98 23 13 98 0.58m
R8 98 23 1.714k
C4 98 23 75f

* 3rd POLE STAGE
G3 98 33 23 98 0.17m
R10 98 33 6k
C5 98 33 75f

* BUFFER STAGE
Gbuf 98 32 33 98 1e-2
Rbuf 98 32 100

* OUTPUT STAGE
R18 25 99 .06
R19 25 50 .06
Vcd 30 25 0
G6 25 99 99 32 16.67
G7 50 25 32 50 16.67
V4 26 25 -.799
V5 25 27 -.799
D5 32 26 Dx
D6 27 32 DX

Fo1 98 70 vcd 1
D7 70 71 DX
D8 72 70 DX
Vi1 98 71 0
Vi2 72 98 0

Erefq 96 0 30 0 1 
Iq 99 50 8.25m
Fq1 99 96 POLY(2) Vi2 Vcd 0 -1 0.5
Fq2 96 50 POLY(2) Vi1 Vcd 0 -1 -0.5

.MODEL QN1 NPN(BF=1000 VA=200 IS=0.5E-15)
.MODEL QN2 NPN(BF=1000 VA=200 IS=0.5E-15)
.MODEL QP1 PNP(BF=1000 VA=200 IS=0.5E-15)
.MODEL QP2 PNP(BF=1000 VA=200 IS=0.5E-15)
.MODEL DX D(IS=1e-15)
.ENDS
