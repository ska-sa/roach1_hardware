*AD8310 SPICE Macro-model
*
*Copyright 2003 by Analog Devices
*
*Refer to "README.DOC" file for License Statement. Use of
*this mod indicates your acceptance of the terms and pro-
*vision in the License Statement.
*
*Node assignments
*		       VPOS
*		       |  INHI
*		       |  |  INLO
*		       |  |  |  COMM
*		       |  |  |  |  ENBL
*		       |  |  |  |  |  BFIN
*		       |  |  |  |  |  |    VOUT
*		       |  |  |  |  |  |    |    OFLT
*		       |  |  |  |  |  |    |    |
*.SUBCKT AD8310 5 1 2 0 7 34 32 80
*Input RC
C1	1	0	1.4p
C2	2	0	1.4p
R1	1	0	1k
R2	2	0	1k
R3	1	13	1E-12
R4	2	13	1E-12
RA	A	0	1k

I_supply	0	8	DC	8mA
R_con_supply	6	8	1E-12
R_supply	5	0	1k

*Slope and Intercept
Vslope 	B 0 .640
Vintercept 	C 0 1.235

*Enable switches
S1	6	5	7	0	ZWIK1
.model ZWIK1 vswitch (RON=1E-12 ROFF=1E12 VON=2V VOFF=0)
S2	A	13	7	0	ZWIK2
.model	ZWIK2	vswitch (RON=1E-12 ROFF=1E12 VON=2V VOFF=0)
V_enable	7	0	2

*Tanh Approximation + Gain Stages
E_TANH1     	41 0 VALUE {0.97*V(B)*TANH(V(C)*(5.188*V(85)))}
E_TANH2     	43 0 VALUE {0.96*V(B)*TANH(V(C)*(5.188*V(42)))}
E_TANH3	45 0 VALUE {0.95*V(B)*TANH(V(C)*(5.188*V(44)))}
E_TANH4	47 0 VALUE {0.99*V(B)*TANH(V(C)*(5.188*V(46)))}
E_TANH5	49 0 VALUE {0.92*V(B)*TANH(V(C)*(5.188*V(48)))}
E_TANH6	51 0 VALUE {1.06*V(B)*TANH(V(C)*(5.188*V(50)))}

E_TANH7	53 0 VALUE {1.70*V(B)*TANH(V(C)*((V(54))))}
E_TANH8	55 0 VALUE {0.198*V(B)*TANH(V(C)*(((V(54))/5.188)))}
E_TANH9	57 0 VALUE {0.21*V(B)*TANH(V(C)*(((V(56))/5.188)))}

*LPF's
R_LPF1	41	42	1k
C_LPF1	42	0	0.01768p
R_LPF2	43	44	1k
C_LPF2	44	0	0.01768p
R_LPF3	45	46	1k
C_LPF3	46	0	0.01768p
R_LPF4	47	48	1k
C_LPF4	48	0	0.01768p
R_LPF5	49	50	1k
C_LPF5	50	0	0.01768p
R_LPF6	51	52	1k
C_LPF6	52	0	0.01768p

R_LPF7	85	54	1k
C_LPF7	54	0	0.01768p
R_LPF8	55	56	1k
C_LPF8	56	0	0.001768p
R_LPF9	57	58	1k
C_LPF9	58	0	0.001768p

*X2
E_X1		71 0 VALUE {(V(42))^2}
E_X2		72 0 VALUE {(V(44))^2}
E_X3		73 0 VALUE {(V(46))^2}
E_X4		74 0 VALUE {(V(48))^2}
E_X5		75 0 VALUE {(V(50))^2}
E_X6		76 0 VALUE {(V(52))^2}

E_X7		77 0 VALUE {0.483*((V(53))^2)}
E_X8		78 0 VALUE {4.95*(V(56))^2}
E_X9		79 0 VALUE {(V(58))^2}

*Offset Compensation Loop
G_loop		80	0	VALUE {V(52)/180k}
C_filt		80	0	20u
R_filt		80	0	16.08154MEG
*R_DC		80	0	1E-6 *Uncomment to allow for DC operation
E_loop		84	0	VALUE {V(80)*(-136/48k)}
E_SUM51	85	0	VALUE	{V(A)+V(84)}

*Summation Functions
E_SUM         	11 0 VALUE {V(71)+V(72)+V(73)+V(74)+V(75)+V(76)+V(77)+V(78)+V(79)}
G_SUM	0 30 VALUE {(V(11)/3k)+.04m}

*Output C/R - LPF
R_R2 		30 0 3k
C_C2		30 0 3p
E_Out		33 0 VALUE {V(30)}
R_Out		33 34 1k
C_Out		34 0   2.768p
Eout1		32 0 VALUE {V(34)}
Rout1		32 0 0.05

VIND 		1 0 sin(0 1 900MEG)
*VIND 		1 0 10

.tran 1n 150n
*.DC DEC VIND 1u 10 500
.OP
.PROBE
.END