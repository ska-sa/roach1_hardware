* AD712J SPICE Macro-model                   4/92, Rev. B
*                                           JCB/JW/PMI
*
* This version of the AD712 model simulates the worst case 
* parameters of the 'J' grade.  The worst case parameters
* used correspond to those in the data sheet.
*
* Revision History:
*     Rev B:  Convert model into ADSpice format
*	         Add noise generators 
*
* Copyright 1990 by Analog Devices, Inc.
*
* Refer to "README.DOC" file for License Statement.  Use of this model
* indicates your acceptance with the terms and provisions in the License Statement.
*
* Node assignments
*                non-inverting input
*                | inverting input
*                | | positive supply
*                | | |  negative supply
*                | | |  |  output
*                | | |  |  |
.SUBCKT AD712J   1 2 99 50 30
*
* INPUT STAGE
*
R3   5  50    5.305
R4   6  50    5.305
CIN  1   2    5.5E-12
I1   99  4    100E-3
IOS  1   2    12.5E-12
EOS  60  1    POLY(1)  17 24  3E-3  1
EN   7  60    42  0  1
GN1  0   1    45  0  1E-6
GN2  0   2    48  0  1E-6
J1   5   2    4   JX
J2   6   7    4   JX
GB1  2  50    POLY(3) 4,2 5,2 50,2 0 1E-12 1E-12 1E-12
GB2  7  50    POLY(3) 4,7 6,7 50,7 0 1E-12 1E-12 1E-12
*
EREF 98  0    24  0   1
*
* VOLTAGE NOISE GENERATOR
*
VN1  41  0    DC 2
DN1  41 42    DEN
DN2  42 43    DEN
VN2  0  43    DC 2
*
* CURRENT NOISE GENERATOR
*
VN3  44  0    DC 2
DN3  44 45    DIN
DN4  45 46    DIN
VN4  0  46    DC 2
*
* CURRENT NOISE GENERATOR
*
VN5  47  0    DC 2
DN5  47 48    DIN
DN6  48 49    DIN
VN6  0  49    DC 2
*  
* SECOND STAGE & POLE AT 32 HZ
*
R5   9  98    7.96E5
C3   9  98    6.25E-9
G1   98  9    5  6  1.88E-1
V2   99  8    2.2
V3   10 50    2.8
D1   9   8    DX
D2   10  9    DX
*
* COMMON-MODE GAIN NETWORK WITH ZERO AT 2.4kHZ
*
R11  16 17     1E6
C8   16 17     6.695E-11
R12  17 98     1
E3   16 98     POLY(2) 1  98  2  98  0  79.24 79.24
*
* POLE AT 15 MHZ
*
R13  18 98     1E3
C9   18 98     10.61E-12
G5   98 18     9  24  1E-3
*
* OUTPUT STAGE
*
R14  24 99     500E3
R15  24 50     500E3
CF   24  0     1E-6
ISY  99 50     -93.2E-3
R16  29 99     110
R17  29 50     110
L1   29 30     1E-8
G6   27 50     18 29  9.09E-3
G7   28 50     29 18  9.09E-3
G8   29 99     99 18  9.09E-3
G9   50 29     18 50  9.09E-3
V4   25 29     0.675
V5   29 26     0.675
D3   18 25     DX
D4   26 18     DX
D5   99 27     DX
D6   99 28     DX
D7   50 27     DY
D8   50 28     DY
F1   29  0     V4  1
F2   0  29     V5  1
*
* MODELS USED
*
.MODEL JX PJF(BETA=1.78E-1  VTO=-2.000  IS=75E-12 RD=0
+ RS=0 CGD=1E-12 CGS=1E-12)
.MODEL DX   D(IS=1E-15 RS=0 CJO=1E-12)
.MODEL DY   D(IS=1E-15 BV=50 RS=10 CJO=1E-12)
.MODEL DEN  D(IS=1E-12 RS=30909 KF=2.651E-15 AF=1)
.MODEL DIN  D(IS=1E-12 RS=12090 KF=0 AF=1)
.ENDS AD712J
