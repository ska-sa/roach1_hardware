*==========================================================
* Analog Devices Linear ICs
*
* This model was developed by:
* AEI Systems, LLC
* 5777 W. Century Blvd. Suite 876
* Los Angeles, California 90045
* Copyright 2002, all rights reserved.
*
* This model is subject to change without notice.
* Users may not directly or indirectly re-sell or 
* re-distribute this model.
*
* For more information contact 
* AEi by email: info@aeng.com. http://www.AENG.com
*
*==========================================================
***************
* |=======================================================
* | ADI LOW NOISE AMPLIFIER MACRO-MODEL AD8331/2/4 LNA
* |=======================================================
*
* Connections:
*
.SUBCKT LNA LMD INH VPSL LON LOP COML COMM ENBL
Q1 1 INH 2 _NPNIN 
I1 VPSL 1 DC=500U
I2 2 COML DC=500U
E1 4 COML 6 1 1MEG
C1 1 LOP1 1.4707P
R1 LOP1 3 0.38889K
V1 VPSL 6 DC=100M
Q2 8 LMD 9 _NPNIN 
I3 VPSL 8 DC=340U
I4 9 COML DC=340U
E2 5 COML 6 8 1MEG
C2 8 LON1 1P
R2 7 LON1 0.5K
VSNSP 2 76 DC=0
F11 COML 78 VSNSP 1
F10 COML 2 VSRP 1
D33 78 79 _DLIM 
VSRP 79 COML DC=4.87
R4 4 LOP1 100
R58 78 COML 10K
R6 76 3 10
E3 CM1 COML VPSL COML 0.5
R8 LMD 10 6K
R3 3 7 0.11111K
R9 INH 10 6K
F13 COML 80 VSNSN 1
I5 COMM VPSL DC=1104.8U
D34 80 81 _DLIM 
VSRN 81 COML DC=3.27
R59 80 COML 10K
R13 25 CM1 1MEG
F12 COML 9 VSRN 1
VSNSN 9 77 DC=0.010167
VSNS1 28 29 DC=0
C8 INH COML 13P
R17 29 LON 5
R5 5 LON1 100
D1 1 VPSL _DLIM 
F1 VPSL 28 VLP1 -1
F2 28 COML VLN1 -1
GB11 CM1 25 Value = {(V(LON1)-V(CM1))*V(ENL1)*1U}
VLN1 0 15 DC=.63
D4 12 14 _DDEF 
D6 14 17 _DDEF 
D5 14 16 _DDEF 
D3 11 14 _DDEF 
R11 13 12 100
R7 7 77 10
R12 15 16 100
VLP1 13 0 DC=.63
V4 17 0 DC=16.36
R15 VPSL LON 100MEG
R16 LON COML 100MEG
R14 25 28 100MEG
V3 0 11 DC=16.36
E7 CM1 COML1 CM1 COML 1
D2 8 VPSL _DLIM 
D11 26 25 _DLIM 
V7 26 COML1 DC=1.34
D12 25 27 _DLIM 
V8 PSL1 27 DC=1.34
V2 10 CM1 DC=0.75
E6 PSL1 CM1 VPSL CM1 1
C9 LMD COML 13P
R22 30 CM1 1MEG
VSNS2 33 34 DC=0
R26 34 LOP 5
F3 VPSL 33 VLP2 -1
F4 33 COML VLN2 -1
GB12 CM1 30 Value = {(V(LOP1)-V(CM1))*V(ENL1)*1U}
VLN2 0 22 DC=.63
D8 19 21 _DDEF 
D10 21 24 _DDEF 
D9 21 23 _DDEF 
D7 18 21 _DDEF 
R20 20 19 100
R21 22 23 100
VLP2 20 0 DC=.63
V6 24 0 DC=16.36
R24 VPSL LOP 100MEG
R25 LOP COML 100MEG
R23 30 33 100MEG
V5 0 18 DC=16.36
D13 31 30 _DLIM 
V9 31 COML1 DC=1.34
D14 30 32 _DLIM 
V10 PSL1 32 DC=1.34
GB9 21 0 Value = {I(VSNS2)*V(ENL1)}
GB10 14 0 Value = {I(VSNS1)*V(ENL1)}
R39 ENBL COML 40K
EB13 74 0 Value = {IF(V(ENBL) - V(COML) < 1.625 , 0 , 1)}
R40 74 ENL1 1K
C6 ENL1 0 10P
G4 VPSL COMM ENL1 0 11M
.MODEL _NPNIN NPN BF=5000 KF=2.5e-14
.MODEL _DDEF D
.MODEL _DLIM D EG=.222 N=.2
.ENDS
