* OP90A SPICE Macro-model                   10/92, Rev. C
*                                           JCB / PMI
*
* Revision History:
*   REV. C
*     Altered gain stage for proper open-loop gain.
*   REV. B
*     Re-ordered subcircuit call out nodes to put the 
*     output node last.
*     Changed Ios from 3E-9 to 1.5E-9
*
*
* This version of the OP-90 model simulates the worst case 
* parameters of the 'A' grade.  The worst case parameters
* used correspond to those in the data book.
*
*
* Copyright 1990 by Analog Devices, Inc.
*
* Refer to "README.DOC" file for License Statement.  Use of this model
* indicates your acceptance with the terms and provisions in the License Statement.
*
* Node assignments
*              non-inverting input
*              | inverting input
*              | | positive supply
*              | | |  negative supply
*              | | |  |  output
*              | | |  |  |
.SUBCKT OP90A  1 2 99 50 31
*
* INPUT STAGE & POLE AT 10 KHZ
*
R1    2  3     5E11
R2    1  3     5E11
R3    5 51     61.6E3
R4    6 51     61.6E3
CIN   1  2     4E-12
C2    5  6     129.2E-12
I1    97 4     1E-6
IOS   1  2     1.5E-9
EOS   9  1     POLY(1)  23 27  150E-6  1
Q1    5  2  7  QX
Q2    6  9  8  QX
R5    7  4     10E3
R6    8  4     10E3
*
EREF  98 0    27  0  1
EPLUS 97 0    99  0  1
ENEG  51 0    50  0  1 
*
* FIRST GAIN STAGE
*
R7   10 98     1E6
G1   98 10     5  6  101.47E-6
D1   10 11     DX
D2   12 10     DX
E1   97 11     POLY(1) 97 27 -1.4 1
E2   12 51     POLY(1) 27 51 -1.4 1
*
* GAIN STAGE & DOMINANT POLE AT 0.323 HZ
*
R8   13 98     2.464E6
C3   13 98     200E-9
G2   98 13     10 27  0.5E-3
H2   97 14     POLY(1) VS2 2.2 -3E3
E5   15 51     POLY(2) (17,51) (97,27) 2.0 1.5 -0.405
D3   13 14     DX
D4   15 13     DX
*
* ZERO-IN ZERO-OUT CLAMP
*
F1   51  17    VS2  -1000
RS1  17  51    1E9
D5   17  51    DX
D6   51  17    DX
*
* NEGATIVE ZERO AT -100 KHZ
*
R9   19 20     1E6
C4   19 20     -1.59E-12
R10  20 98     1
E3   19 98     13 27  1E6
*
* ZERO - POLE PAIR AT 28 KHZ / 100 KHZ
*
R11  21 22     1E6
L1   22 98     4.09
R12  22 98     2.57E6
G3   98 21     20 27  1E-6
*
* COMMON-MODE GAIN NETWORK WITH ZERO AT 126 HZ
*
R13  23 24     1E6
L2   24 98     1.257E3
G4   98 23     3  27  1E-11
D8   23 97     DX
D9   51 23     DX
*
* ZERO - POLE PAIR AT 40 KHZ / 160 KHZ
*
R14  25 26     1E6
L3   26 98     2.98
R15  26 98     3E6
G5   98 25     21 27  1E-6
*
* OUTPUT STAGE
*
ISY  99 50     8.444E-6
R16  27 99     2.7E6
R17  27 50     2.7E6
R18  30 99     6000
R19  30 50     6000
VS2  30 31     DC 0
G6   28 50     25 30  166.7E-6
G7   29 50     30 25  166.7E-6
G8   30 99     99 25  166.7E-6
G9   50 30     25 50  166.7E-6
D10  99 28     DX
D11  99 29     DX
D12  50 28     DY
D13  50 29     DY
*
* MODELS USED
*
.MODEL QX PNP(BF=33.333)
.MODEL DX   D(IS=1E-15)
.MODEL DY   D(IS=1E-15 BV=50)
.ENDS
