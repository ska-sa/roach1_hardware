.SUBCKT AD8045    1   2   81   101  102  
*                IN+  IN- OUT  VCC  VEE
*
***************************************
* Analog Devices AD8045
* 2004.10.8 v2
* OP AMP modeling services provided by:
* Interface Technologies
* www.i-t.com
***************************************
*
* CMR INPUT
RCM15	1	105	10MEG
RCM25	2	105	10MEG
EOS	1 92	POLY(1) 300 100	  0 1
Q1	5 9	7	NPN
Q2	6 2	8	NPN
RC1	101	5	537.15 T_ABS=-250
RC2	101	6	537.15
RE1	7	4	485.45
RE2	8	4	485.45
I1	4	102	0.001
Cpeek 2 0 0.5pf
*
* OPEN-LOOP GAIN, FIRST POLE (252KHz) AND SLEW RATE (1350V/u)
G1	100 10	6 5 0.001861684
RP1	10	100	7.585e5
CP1	10	100	7.40741e-7u
*
* CLIPPING OF VOLTAGE OUTPUTS TO RAILS
DP	10 	103	DLIM
VP	101	103	DC	1.654
DN	104	10	DLIM
VN	104	102	DC	1.654
.MODEL DLIM D(IS=1E-15)
*
* NOISE
EN   92 9     36  0  2
GN1  0  2     94  0  .02
GN2  0  1     97  0  .02
*
* VOLTAGE NOISE SOURCE
*
DN1  35 36    DEN
DN2  36 37    DEN
VN1  35  0    DC 2
VN2  0  37    DC 2
*
* CURRENT NOISE SOURCE 1
*
DN3  93 94    DIN
DN4  94 95    DIN
VN3  93  0    DC 2
VN4  0  95    DC 2
*
* CURRENT NOISE SOURCE 2
*
DN5  96 97    DIN
DN6  97 98    DIN
VN5  96  0    DC 2
VN6  0  98    DC 2
*
.MODEL DEN  D(IS=1E-12 RS=5e0 KF=5E-11 AF=1)
.MODEL DIN  D(IS=1E-12 RS=.5e0 KF=0.7e-12 AF=1)
*
*
* COMMON MODE REJECTION GAIN AND POLE: 2Mhz
GCM22	100 300	105 100 5.01E-7
RCM22	300	301	1e2
LCM22	301	100	7.9577E-6
*
*
* 2ND POLE 1.1ghz
G2	100 40	10 100 0.01
RP2	40	100	100
CP2	40	100	1.4469e-12
*
* SUPPLY CURRENT CORRECTION
D1	101	15	DNOM
GSC1	15 100	80 81	0.02
DZ11	100	15	DZ
RZ11    100     15      1MEG
GSC2	100 16	80 81	-0.02
DZ12	16	100	DZ
RZ12    16      100     1MEG
D2	16	102	DNOM
*
.MODEL	DNOM	D(IS=1E-15)
.MODEL	DZ	D(IS=1E-15 BV=50)
*
* CURRENT LIMITING OF OUTPUT
DL1	40	82	DILIM		; 40 IS THE STAGE BEFORE THE OUPUT
VL1	82	81	DC	7.736V 	; 81 IS THE OUPUT PIN, AFTER rOUT
DL2	83	40	DILIM	
VL2	81	83	DC	7.736v
.MODEL 	DILIM	D(IS=1E-15)
*
* OUTPUT STAGE
EOUT	80 100	40 100	1
RO	80	81	50
*
* INTERNAL REFERENCE
RREF1	101	103	100K
RREF2	103	102	100K
EREF	100 0	103 0 1
R100	100	0	1MEG
*
.model NPN  NPN(BF=250)
*
.ENDS
