* SSM2275 SPICE Macro-Model Typcial Values
* 8/97, Ver. 1
* TAM / ADSC
*
* Node assignments
*		noninverting input
*		|	inverting input
*		|	|	positive supply
*		|	|	|	negative supply
*		|	|	|	|	output
*		|	|	|	|	|
*		|	|	|	|	|
.SUBCKT SSM2275 1	2	99	50	45
*
* INPUT STAGE
*
Q1  4  3  5 QNIX
Q2  6  2  7 QNIX
RC1   99 11 15E3
RC2   99 12 15E3
RE1    5  8 1E3
RE2    7  8 1E3
EOS    3  1 POLY(2) (61,98) (73,98) 1E-3 1.78E-5 1
IOS    1  2 5E-9
ECMH1  4 11 POLY(1) (99,50) 0.9 -30E-3
ECMH2  6 12 POLY(1) (99,50) 0.9 -30E-3
ECML1  9 50 POLY(1) (99,50) 0.1 30E-3
ECML2 10 50 POLY(1) (99,50) 0.1 30E-3
D1     9  5 DX
D2    10  7 DX
D3    13  1 DZ
D4     2 13 DZ
IBIAS  8 50 200E-6
*
* CMRR=115 dB, ZERO AT 1kHz, POLE AT 10kHz
*
ECM1 60 98 POLY(2) (1,98) (2,98) 0 .5 .5
RCM1 60 61 159.2E3
RCM2 61 98 17.66E3
CCM1 60 61 1E-9
*
* PSRR=120dB, ZERO AT 400Hz
*
RPS1 70  0 1E6
RPS2 71  0 1E6
CPS1 99 70 1E-5
CPS2 50 71 1E-5
EPSY 98 72 POLY(2) (70,0) (0,71) 0 1 1
RPS3 72 73 1.59E6
CPS3 72 73 250E-12
RPS4 73 98 1.59
*
* INTERNAL VOLTAGE REFERENCE
*
RSY1 99 91 100E3
RSY2 50 90 100E3
VSN1 91 90 DC 0
EREF 98  0 (90,0) 1
GSY  99 50 POLY(1) (99,50) 0.97E-3 -7E-6
*
* ADAPTIVE POLE AND GAIN STAGE
* AT Vsy= 5, fp=12.50MHz,Av=1
* AT Vsy=30, fp=18.75MHz,Av=1.16
*
G2  98 20 POLY(2) (4,6) (99,50) 0 80.3E-6 0 0 2.79E-6
VR1 20 21 DC 0
H1  21 98 POLY(2) VR1 VSN1 0 11.317E3 0 0 -28.29E6
C2  20 98 1.2E-12
*
* POLE AT 90MHz
*
G3 98 23 (20,98) 565.5E-6
R5 23 98 1.768E3
C3 23 98 1E-12
*
* GAIN STAGE
*
G1 98 30 (23,98) 733.3E-6
R1 30 98 9.993E3
CF 30 45 200E-12
D5 31 99 DX
D6 50 32 DX
V1 31 30 0.6
V2 30 32 0.6
*
* OUTPUT STAGE
*
Q3  46 42 99 QPOX
Q4  47 44 50 QNOX
RO1 46 48 30
RO2 47 49 30
VO1 45 48 15E-3
VO2 49 45 10E-3
RB1 41 42 200
RB2 43 44 200
EO1 99 41 POLY(1) (98,30) 0.7528 1
EO2 43 50 POLY(1) (30,98) 0.7528 1
*
* MODELS
*
.MODEL QNIX NPN(IS=1E-16,BF=400,KF=1.96E-14,AF=1)
.MODEL QNOX NPN(IS=1E-16,BF=100,VAF=130)
.MODEL QPOX PNP(IS=1E-16,BF=100,VAF=130)
.MODEL DX D(IS=1E-16)
.MODEL DZ D(IS=1E-14,BV=6.6)
.ENDS SSM2275