* REF02C SPICE MACROMODEL                    9/91, Rev. A
*                                            (JCB / PMI)    
*
* This version of the REF02 model simulates the worst case 
* parameters of the 'C' grade.  The worst case parameters
* used correspond to those in the data sheet.
*
* Copyright 1991 by Analog Devices, Inc.
*
* Refer to "README.DOC" file for License Statement.  Use of this model
* indicates your acceptance with the terms and provisions in the License Statement.
*
*  NODE NUMBERS
*               VIN
*               |  GND
*               |  |  TRIM
*               |  |  |  VOUT
*               |  |  |  |
.SUBCKT REF02C  2  4  5  6
*
* 1.23V REFERENCE
*
I1     4  10   3.6095E-7
R1     10  4   3400E3  TC=65E-6
G1     4  10   21  4  1E-6
F1     4  10   VS  54.6E-9
*
* LINE REGULATION ZERO
*
E1     20  4   2  4  54.6
R11    20 21   1E6
R12    21  4   1
C4     20 21   27E-8
*
* INTERNAL OP AMP
*
G2     4  11   10  19  2E-3
R2     4  11   150E6
C1     4  11   2.6E-10
D1     11 12   DX
V1     2  12   1.9
*
* SECONDARY POLE
*
G3     4  13   11  4  1E-6
R3     4  13   1E6
C2     4  13   2.4E-13
*
* OUTPUT STAGE
*
ISY    2   4   0.985E-3
FSY    2   4   V1  -1 
G4     4  14   13  4  25E-6
R4     4  14   40E3
R7     17 19   6.0488E3
R8     19  4   2E3
R9     19  5   56.0E3
R10    5   4   1E12
Q1     16 14   17   QN
VS     18 17   DC 0
L1     18  6   1E-7
*
* OUTPUT CURRENT LIMIT
*
Q2     15  2   16  QN
R6     2  16   19
R5     2  15   18E3
C3     2  15   1E-6
G5     14  4   2  15  1
*
.MODEL  QN  NPN(IS=1E-15  BF=1000)
.MODEL  DX  D(IS=1E-18)
.ENDS
