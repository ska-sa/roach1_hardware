*****************
* This model was developed for Analog Devices by:
* AEI Systems, LLC
* 5777 W. Century Blvd., Suite 876
* Los Angeles, California  90045-5677
*
* The model is �2006, AEi Systems, LLC. All rights reserved. 
*
* Users may not directly or indirectly display, re-sell or 
* re-distribute this model or any derivative work therefore 
* without the prior written consent of both AEi Systems and 
* Analog Devices. This model is subject to change without 
* notice. Neither Analog Devices nor AEi Systems is responsible 
* for updating this model.
*
* For more information regarding modeling services, model 
* libraries and simulation products, please call AEi Systems 
* at (310) 216-1144, or contact AEi Systems by 
* email: info@aeng.com. Or visit AEi Systems on the web 
* at http://www.AENG.com


*$
.SUBCKT AD737 CC VIN PD NVS COM VS VOUT CAV

* Use .OPTIONS GMIN=5E-17 for best output accuracy

R1 3 13 8K
R3 3 1 4K
R4 1 15 3K
Q1 VS 4 15 NPN
.MODEL NPN NPN
R9 6 13 3K
ER VOUT II Value={IF(V(PD) < V(VS), 1U*I(VER), 1G*I(VER))}
VER II 16
GB3 COM CAV Value={I(V4)*I(V4)}
R5 10 NVS 8K
V5 CAV 10
GB1 16 COM Value={IF(V(PD) < V(VS), (IF(SQRT(I(V5)) > 1.7/8000, 1.7/8000, SQRT(I(V5)))), 0)}
R6 CC 18 8K
RPD PD 0 1G
X2 1 COM 4 VS NVS AEIOPAMP0 
Q7 VS 4 6 NPN
V4 13 COM
R10 16 COM 8K
GB2 0 VIN VALUE={1P + 50P*V(VIN)}
GB4 0 18 VALUE={1P + 5P*V(CC)}
EB5 3 0 VALUE={IF(ABS(V(VIN)) > ABS(V(CC)), V(VIN), V(CC))}
.ENDS
*$
.SUBCKT AEIOPAMP0 2    3  6   7   4
RP 4 7 10K
IB 3 90 5.0000N
VIB 90 4
IO 3 2 500.00P
RIP 3 4 1G
CIP 3 4 1.4PF
FIBN 2 4 VIB 1
RIN 2 4 1G
CIN 2 4 1.4PF
VOFST 2 10 10.0000N
RID 10 3 1G
EA 11 4 10 3 1
R1 11 12 5K
R2 12 13 50K
C1 12 4 130.00F
GA 4 14 4 13 202.50 
C2 13 14 27.000F
RO 14 4A 75
EBAL 4A 4 2A 4 1
RBAL1 7 2A 1MEG
RBAL2 2A 4 1MEG
L 14 6 300.00N
RL 14 6 1000
CL 6 4 3PF
D1 6 70 DN
VSAT 70 7 -1.0000 
D2 40 6 DN
VSAT2 40 4 3.0000 
.MODEL DN D
.ENDS
*$

