* OP467G SPICE Macro-model             5/92, Rev. A
*                                       ARG / PMI
*
* Copyright 1993 by Analog Devices
*
* Refer to "README.DOC" file for License Statement.  Use of
* this model indicates your acceptance of the terms and pro-
* visions in the License Statement.
*
* Node assignments
*                non-inverting input
*                |  inverting input
*                |  |  positive supply
*                |  |  |  negative supply
*                |  |  |  |  output
*                |  |  |  |  |
.SUBCKT OP467G   1  2  99 50 27
*
* INPUT STAGE
*
I1   4    50   10E-3
CIN  1    2    1E-12
IOS  1    2    50E-9
Q1   5    2    8    QN
Q2   6    7    9    QN
R3   99   5    66.472
R4   99   6    66.472
R5   8    4    61.3
R6   9    4    61.3
EOS  7    1    POLY(1) (14,20) 0.5E-3 4
EREF 98   0    (20,0) 1
*
* GAIN STAGE AND DOMINANT POLE AT 2.12KHZ
*
R7   10   0    938.942E3
C2   10   0    80E-12
G1   0    10   (5,6) 15.044E-3
V1   99   11   2.025
V2   12   50   2.025
D1   10   11   DX
D2   12   10   DX
RC   10   28   1.4E3
CC   28   27   12E-12
*
* COMMON MODE STAGE WITH ZERO AT 5.024KHZ
*
ECM  13   98   POLY(2) (1,20) (2,20) 0 0.5 0.5
R8   13   14   1E6
R9   14   98   25.119
C3   13   14   31.680E-12
*
* POLE AT 400E6
*
R10  15   98   1E6
C4   15   98   0.398E-15
G2   98   15   (10,20) 1E-6
*
* OUTPUT STAGE
*
ISY  99   50   -7.656E-3
RMP1 99   20   96.429E3
RMP2 20   50   96.429E3
RO1  99   26   200
RO2  26   50   200
L1   26   27   1E-7
GO1  26   99   (99,15) 5E-3
GO2  50   26   (15,50) 5E-3
G4   23   50   (15,26) 5E-3
G5   24   50   (26,15) 5E-3
D5   99   23   DX
D6   99   24   DX
D7   50   23   DY
D8   50   24   DY
*
* MODELS USED
*
.MODEL QN NPN(BF=8.333E3)
.MODEL DX D
.MODEL DY D(BV=50)
.ENDS
