*ADG513_5 Spice Macromodel                        5/95
*                                              WF/ADSC
*
*  This Macromodel should be used for simulating the operation
*  of the ADG513 with a single +5 Volt power supply.
*     For Single +3 V operation, use the ADG513_3.CIR Macromodel
*     For �5 V operation, use the ADG513�5.CIR Macromodel
*     For �15 V operation, use the ADG413.CIR Macromodel
*
*
* Copyright 1995 by Analog Devices, Inc.
*
* Refer to "README.DOC" file for License Statement.
* Use of this model indicates your acceptance of
* the terms and provisions in the License Statement.
*
* Node assignments
*                  IN1 
*                  | D1
*                  | | S1
*                  | | | VSS
*                  | | | | GND
*                  | | | | | S4
*                  | | | | | | D4
*                  | | | | | | | IN4
*                  | | | | | | | | IN3
*                  | | | | | | | | | D3
*                  | | | | | | | | | |  S3
*                  | | | | | | | | | |  |  VL
*                  | | | | | | | | | |  |  |  VDD
*                  | | | | | | | | | |  |  |  |  S2
*                  | | | | | | | | | |  |  |  |  |  D2
*                  | | | | | | | | | |  |  |  |  |  |  IN2
*                  | | | | | | | | | |  |  |  |  |  |  |
.SUBCKT ADG513_5   1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
*
* SWITCH 1
*
MP1   20  1   12  12  PCNTRL  L=6E-6 W=90E-6
MN1   20  1   5   5   NCNTRL  L=6E-6 W=210E-6
IL1   1   5   5E-9
C1    20  4   120P
MP2   21  22  13  13  PCNTRL  L=6E-6 W=20E-6
MN2   21  22  4   4   NCNTRL  L=6E-6 W=20E-6
C2    21  4   20P
E1    22  26  POLY(2) (20,5) (12,5) 0 9 -4.5
E2    26  0   POLY(2) (13,0) (4,0) 0 0.5 0.5
MP3   2   24  3   13   PSW  L=6E-6 W=1600E-6
MN3   2   25  3   4    NSW  L=6E-6 W=3038E-6
EPN1  24  13  21  4   -1
ECN1  25  13  13  21  -1
CS1   3   5   7.4E-12
CD1   2   5   7.4E-12
CSD1  2   3   1.3E-12
*
* SWITCH 2
*
MP4   30  16  12  12  PCNTRL  L=6E-6 W=90E-6
MN4   30  16  5   5   NCNTRL  L=6E-6 W=210E-6
IL2   16  5   5E-9
C3    30  4   120P
MP5   31  32  13  13  PCNTRL  L=6E-6 W=20E-6
MN5   31  32  4   4   NCNTRL  L=6E-6 W=20E-6
C4    31  4   20P
E3    32  36  POLY(2) (30,5) (12,5) 0 9 -4.5
E4    36  0   POLY(2) (13,0) (4,0) 0 0.5 0.5
MP6   15  34  14  13   PSW  L=6E-6 W=2000E-6
MN6   15  35  14  4    NSW  L=6E-6 W=1000E-6
EPN2  34  4   31  4   1
ECN2  35  4   13  31  1
CS2   14  5   7.4E-12
CD2   15  5   7.4E-12
CSD2  15  14  1.3E-12
*
* SWITCH 3
*
MP7   40  9   12  12  PCNTRL  L=6E-6 W=90E-6
MN7   40  9   5   5   NCNTRL  L=6E-6 W=210E-6
IL3   9   5   5E-9
C5    40  4   120P
MP8   41  42  13  13  PCNTRL  L=6E-6 W=20E-6
MN8   41  42  4   4   NCNTRL  L=6E-6 W=20E-6
C6    41  4   20P
E5    42  46  POLY(2) (40,5) (12,5) 0 9 -4.5
E6    46  0   POLY(2) (13,0) (4,0) 0 0.5 0.5
MP9   10  44  11  13   PSW  L=6E-6 W=2000E-6
MN9   10  45  11  4    NSW  L=6E-6 W=1000E-6
EPN3  44  4   41  4   1
ECN3  45  4   13  41  1
CS3   11  5   7.4E-12
CD3   10  5   7.4E-12
CSD3  10  11  1.3E-12
*
* SWITCH 4
*
MP10  50  8   12  12  PCNTRL  L=6E-6 W=90E-6
MN10  50  8   5   5   NCNTRL  L=6E-6 W=210E-6
IL4   8   5   5E-9
C7    50  4   120P
MP11  51  52  13  13  PCNTRL  L=6E-6 W=20E-6
MN11  51  52  4   4   NCNTRL  L=6E-6 W=20E-6
C8    51  4   20P
E7    52  56  POLY(2) (50,5) (12,5) 0 9 -4.5
E8    56  0   POLY(2) (13,0) (4,0) 0 0.5 0.5
MP12  7   54  6   13   PSW  L=6E-6 W=2000E-6
MN12  7   55  6   4    NSW  L=6E-6 W=1000E-6
EPN4  54  13  51  4   -1
ECN4  55  13  13  51  -1
CS4   6   5   7.4E-12
CD4   7   5   7.4E-12
CSD4  7   6   1.3E-12
*
* CROSSTALK CAPACITORS
CS12  3   14   0.12E-12
CD12  2   15   0.12E-12
CS13  3   11   0.12E-12
CD13  2   10   0.12E-12
CS14  3   6    0.12E-12
CD14  2   7    0.12E-12
CS23  14  11   0.12E-12
CD23  15  10   0.12E-12
CS24  14  6    0.12E-12
CD24  15  7    0.12E-12
CS34  11  6    0.12E-12
CD34  10  7    0.12E-12
*
.MODEL  PCNTRL  PMOS(VTO=-1 RD=0.1 RS=0.1)
.MODEL  NCNTRL  NMOS(VTO=1 RD=.1 RS=.1)
.MODEL  PSW     PMOS(LEVEL=1 VTO=-.5 GAMMA=0.3772 PHI=0.5 RS=5
+ UO=279.4 TOX=100E-9 LAMBDA=0.3141 CGSO=172.6E-12 kp=4.5E-5
+ CGDO=172.6E-12 CGBO=69.1E-12 CJ=120E-12
+ CJSW=597E-6 JS=3.2E-6 KF=1E-30 AF=1)
.MODEL  NSW     NMOS(LEVEL=1 VTO=.3 GAMMA=1.412 PHI=0.7 RS=15
+ UO=662.6 TOX=100E-9 LAMBDA=.013 CGSO=172.6E-12 KP=3.5E-5
+ CGDO=172.6E-12 CGBO=69.1E-12 CJ=170E-6
+ CJSW=298E-6 JS=2.7E-6 KF=3.6E-29 AF=1)
.ENDS ADG513_5
.END
