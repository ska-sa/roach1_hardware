* AD8033 Spice Model		Rev. 0	VC
* Refer to "README.DOC" file for License Statement.
* Use of this model indicates your acceptance with
* the terms and provisions in the License Statement.
*
* The following parameters are accurately modeled;
*
*       closed loop gain vs. frequency
*       output clamping voltage and current
*	     input common mode range for FET input
*       input impedance
*       slew rate
*       output currents are reflected to V supplies
*       Vos is static and will not vary
*       Ibias current will remain around 50 pA over common mode range
*       distortion is not characterized       
*
*
*
*    Node assignments
*              non-inverting input
*              | inverting input
*              | | positive supply
*              | | |  negative supply
*              | | |  |  output
*              | | |  |  |
.SUBCKT AD8033 1 2 99 50 30
				 
* FET INPUT STAGE


Vos 9 2 1e-3
Ios 2 1 0.75e-6
Cd 1 2 1.7p
Ccm1 1 0 2.3p
Ccm2 2 0 2.3p
J1 5 1 10 NMOD 
J2 6 9 11 NMOD 
R3 99 5 1132 
R4 99 6 1132
R5 10 4 1020
R6 11 4 1020
I11 4 50 225u
			  
* GAIN STAGE & POLE AT 2.47 kHz
Eref 15 0 POLY(2) 99 0 50 0 0 .5 .5 
G1 13 15 5 6 1
R7 13 15 28k
C3 13 15 2.3n
V1 98 14 0.12
V2 16 52 0.12
D1 13 14 DX
D2 16 13 DX

Ecc 98 0 99 0 1
Ess 52 0 50 0 1

*POLE AT 350 MHz
G2 15 43 13 15 440e-6
R10 15 43 2.27k
C5 15 43 0.2p

*POLE AT 425 MHz
G3 15 53 43 15 534e-6
R11 15 53 1.87k
C6 15 53 0.2p

*POLE AT 834 MHz
G4 15 63 13 15 628e-6
R12 15 63 1.59k
C7 15 63 0.12p

* BUFFER STAGE
Gbuf 15 32 63 15 1e-3
Rbuf 32 15 1000

* OUTPUT STAGE
Vo1 99 90 0
Vo2 51 50 0
R18 25 90 .04
R19 25 51 .04
Vcd 25 30 0
G6 25 90 99 32 25
G7 51 25 32 50 25
V4 26 25 -0.846
V5 25 27 -0.846
D5 32 26 Dx
D6 27 32 DX

Fo1 15 70 vcd 1
D7 70 71 DX
D8 72 70 DX
Vi1 71 15 0
Vi2 15 72 0

Erefq 96 0 30 0 1 
Iq 99 50 3.08m
Fq1 96 99 POLY(2) Vo1 Vi1 0 1 -1
Fq2 50 96 POLY(2) Vo2 Vi2 0 1 -1

.MODEL NMOD NJF VTO=0.222 BETA=100 IS=1e-14
.MODEL DX D(IS=1e-15) 
.ENDS
