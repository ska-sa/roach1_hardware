* AD824 SPICE Macro-model               9/94, Rev. A
*                                       ARG / PMI
*
* Copyright 1993 by Analog Devices, Inc.
*
* Refer to "README.DOC" file for License Statement.  
* Use of this model indicates your acceptance with 
* the terms and provisions in the License Statement.
*
* Node assignments
*                non-inverting input
*                |  inverting input
*                |  |  positive supply
*                |  |  |  negative supply
*                |  |  |  |  output
*                |  |  |  |  |
.SUBCKT AD824    1  2  99 50 25
*
* INPUT STAGE & POLE AT 3.1MHZ
*
R3   5    99   1.193E3
R4   6    99   1.193E3
CIN  1    2    4E-12
C2   5    6    19.229E-12
I1   4    50   108E-6
IOS  1    2    1E-12
EOS  7    1    POLY(1) (12,98) 100E-6 1
J1   4    2    5    JX
J2   4    7    6    JX
*
* GAIN STAGE & DOMINANT POLE
*
EREF 98   0    (30,0) 1
R5   9    98   2.205E6
C3   9    25   54E-12
G1   98   9    (6,5) 0.838E-3
V1   8    98   -1
V2   98   10   -1
D1   9    10   DX
D2   8    9    DX
*
* COMMON-MODE GAIN NETWORK WITH ZERO AT 1KHZ
*
R21  11   12   1E6
R22  12   98   100
C14  11   12   159E-12
E13  11   98   POLY(2) (2,98) (1,98) 0 0.5 0.5
*
* POLE AT 10MHZ
*
R23  18   98   1E6
C15  18   98   15.9E-15
G15  98   18   (9,98) 1E-6
*
* OUTPUT STAGE
*
ES   26   98   (18,98) 1
RS   26   22   500
IB1  98   21   2.404E-3
IB2  23   98   2.404E-3
D10  21   98   DY
D11  98   23   DY
C16  20   25   2E-12
C17  24   25   2E-12
DQ1  97   20   DQ
Q2   20   21   22  NPN
Q3   24   23   22  PNP
DQ2  24   51   DQ
Q5   25   20   97  PNP 20
Q6   25   24   51  NPN 20
VP   96   97   0
VN   51   52   0
EP   96   0    (99,0) 1
EN   52   0    (50,0) 1
R25  30   99   5E6
R26  30   50   5E6
FSY1 99   0    VP 1
FSY2 0    50   VN 1
DC1  25   99   DX
DC2  50   25   DX
*
* MODELS USED
*
.MODEL JX NJF(BETA=3.2526E-3 VTO=-2.000 IS=2E-12)
.MODEL NPN NPN(BF=120 VAF=150 VAR=15 RB=2E3
+ RE=4 RC=550 IS=1E-16)
.MODEL PNP PNP(BF=120 VAF=150 VAR=15 RB=2E3
+ RE=4 RC=750 IS=1E-16)
.MODEL DX D(IS=1E-15)
.MODEL DY D()
.MODEL DQ D(IS=1E-16)
.ENDS AD824
