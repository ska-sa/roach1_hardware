*  AD8016 Spice Macro-model                  DATE JUNE 27,00  
* Rev A
*															JCH, ADI Cent Apps
*  Copyright 1998 by Analog Devices, Inc.
*
* Refer to "README.DOC" file for License Statement.
* Use of this model indicates your acceptance with
* the terms and provisions in the License Statement.
*
*CAUTION: Pwrdn0 AND Pwrdn1 ARE DIGITAL CONTROLS FOR
*REDUCING POWER CONSUMPTION.  EXERCISING THESE 
*CONTROLS HAS NO EFFECT ON FREQUENCY RESPONSE.
*
* Node assignments
*                non-inverting input
*                | inverting input
*                | | positive supply
*                | | |  negative supply
*                | | |  |  output
*                | | |  |  |  Pwrdn0
*                | | |  |  |  | Pwrdn1
*                | | |  |  |  | |
.SUBCKT AD8016t5  1 2 99 50 61 5 6


***** Input Stage

q1 4 4 41 qn1 
q2 3 3 41 qp1
i1 99 4 3e-4
i2 3 50 3e-4

*cin1 4 88 1.5pf
*cin2 2 88 1.5pf

q3 9 4 2 qn2
q4 10 3 2 qp2

rxxa 99 4 100k
rxxb 3 50 100k
  

VT1  9  99 0   
VT2 10 50 0  

vos 41 1 0
*eos 41 1 poly(1) 43 88 5e-3 1

***** internal vnoise source

*dn1 42 88 dnv
*rn1 42 88 5e-3
*vn1 42 88 0

*hn1 43 88 vn1 1
*rn2 43 88 1

***** internal inoise source

*dn2 72 88 dniinv
*rn3 72 88 50
*vn2 72 88 0

*hn2 73 88 vn2 1
*rn4 73 88 1

***** internal reference

Eref 88 0 poly(2) 99 0 50 0 0 0.5 0.5

***** gain stage/dominant pole/clamp circuitry

F3 29 88 VT1 1 
F4 29 88 VT2 1  
r3 29 88 1meg
c1 29 88 8.03f

vc1 99 45 1.33
vc2 46 50 1.31
dc1 29 45 dx
dc2 46 29 dx

***** pole at 114MHz

egain2 32 88 88 29 1
r4 32 44 1
c3 44 88 1.2n

***** pole at 114MHz

*egain3 33 88 32 88 1
*r5 33 47 1
*c4 47 88 1.4n

***** buffer to output stage

gbuf 34 88 44 88 1e-2
re1 34 88 100

*****output current mirroring to supplies

fo1 88 110 vcd 1
do1 110 111 dx
do2 112 110 dx
vi1 111 88 0
vi2 88 112 0
fsy1 99 0 poly(2) visy1 vi1 0 -1 1
fsy2 0 50 poly(2) visy2 vi2 0 -1 1
isy1 99 0 2.84m
isy2 0 50 3.08m

S1 99 36 6 0 SW13
S2 36 0 6 0 SW24
Isw1  36 0 2.55m

S3 99 37 5 0 SW13
S4 37 0 5 0 SW24
Isw2 37 0 5.55m

S5 50 38 6 0 SW13
S6 38 0 6 0 SW24
Isw3 0 38 2.5m

S7 50 39 5 0 SW13
S8 39 0 5 0 SW24
Isw4 0 39 5.5m

Rlog1 99 5 100k
Rlog2   5 0 100k
Rlog3 99 6 100k
Rlog4   6 0 100k


***** output stage

go3 60 63 99 34 0.385
go4 64 60 34 50 0.385
r03 60 63 2.6 
r04 60 64 2.6 
visy1 99 63 0
visy2 64 50 0
vcd 60 61 0   
*lo1 62 61 1e-10
do5 34 70 dx
do6 71 34 dx
vo1 70 60 -0.083
vo2 60 71 -0.085

.model dx d(is=1e-13 kf=1e-30)
.model dy d(is=26e-9 kf=1e-30)
.model dnv d(is=1e-15 kf=2e-15 af=0)
.model dniinv d(is=1e-15 kf=1e-19 af=0)
.model qn1 npn(bf=200 kf=1e-30 af=0)
.model qn2 npn(bf=200 kf=1e-30 af=0)
.model qp1 pnp(bf=200 kf=1e-30 af=0)
.model qp2 pnp(bf=200 kf=1e-30 af=0)
.model SW13 vswitch ron=0.1 roff=1meg von=1.6 voff=1.5
.model SW24 vswitch ron=100 roff=1meg von=1.5 voff=1.6
.ends ad8016t5
