* AD584L SPICE Macromodel 1/2001, Rev. B
* AAG / PMI
* TRW / PMI
*
* This version of the AD584 voltage reference model simulates the worst case
* parameters of the 'L' grade.  The worst case parameters used correspond
* to those parameters in the data sheet.
*
* Copyright 1993 by Analog Devices, Inc.
*
* Refer to "README.DOC" file for License Statement.  Use of this model
* indicates your acceptance with the terms and provisions in the License Statement.
*
*  NODE NUMBERS
*              10.0 V
*              |  5.0 V
*              |  |  2.5 V
*              |  |  |  GND
*              |  |  |  |  STROBE
*              |  |  |  |  |  VBG
*              |  |  |  |  |  |  CAP
*              |  |  |  |  |  |  |  VIN
*              |  |  |  |  |  |  |  |
.SUBCKT AD584L 1  2  3  4  5  6  7  8
*
* BANDGAP REFERENCE
*
I1 4 10 DC 1.214243E-3
R1 10 4 1E3 TC=5E-6
EN 10 11 41 0 1
G1 4 11 8 4 2.430243E-8
F1 4 11 POLY(2) VS1 VS2 (0,6.0756E-5,6.0756E-5)
*
* NOISE VOLTAGE GENERATOR
*
VN1 40 0 DC 2
DN1 40 41 DEN
CN 41 0 50E-12
DN2 41 42 DEN
VN2 0 42 DC 2
*
* INTERNAL OP AMP AND DOMINANT POLE @ 5 Hz
*
G2 4 7 11 6 1E-3
R2 7 4 1E8
C1 7 4 3.1831E-10
D1 7 12 DX
V1 8 12 DC 1.5
*
* SECONDARY POLE @ 1 MHz
*
G3 4 13 7 4 1E-6
R3 13 4 1E6
C2 13 4 1.5915E-13
*
* OUTPUT STAGE
*
ISY 8 4 6.015E-4
FSY 8 4 V1 -1
*
G4 4 14 13 4 20E-6
R4 14 4 50E3
FSC 14 4 VSC 1
Q1 4 14 5 QP
I2 8 5 DC 100E-6
VSC 8 15 DC 0
QSC 15 8 16 QN
RSC 8 16 24.5
Q2 16 5 17 QN
VS1 19 17 DC 0
Q3 4 5 18 QP
VS2 18 19 DC 0
R5 19 2 25.0005k
R6 2 3 12.49995k
R7 3 6 6.42405k
R8 6 4 6.075k
LO 19 1 1E-7
*
.MODEL QN NPN(IS=1E-15 BF=1E3)
.MODEL QP PNP(IS=1E-15 BF=1E3)
.MODEL DX D(IS=1E-15)
.MODEL DEN D(IS=1E-12 RS=4.56436E5 AF=1 KF=2.81234E-17)
.ENDS AD584L
