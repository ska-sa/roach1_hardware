* OP2177 SPICE Macro-model              
*  05/02 Rev A
* SB, ADSiV apps                                    
* Typical values, Vsy=�15V
* Copyright 2002 by Analog Devices
*
* Refer to "README.DOC" file for License Statement.  Use of this model
* indicates your acceptance with the terms and provisions in the License Statement.
*
* Node assignments
*               non-inverting input
*               | inverting input
*               | | positive supply
*               | | |  negative supply
*               | | |  |  output
*               | | |  |  |
*               | | |  |  |
.SUBCKT OP2177  1 2 99 50 34
*
* INPUT STAGE & POLE AT 100 MHZ
*
R3   5 51     6.8E3
R4   6 51     6.8E3
CIN  1  2     1.5E-12
C2   5  6      3.5E-12
I1   97 4      500E-6
IOS  1  2     0.1E-9
EOS  9  3     POLY(2)  (26, 28) (73, 98) 15E-6  1 1
Q1   5  2  7  QX
Q2   6  9  8  QX
R5   7  4     50
R6   8  4     50
D1   2 36     DZ
D2   1 36     DZ
EN   3  1     10  0  1
GN1  0  2     13  0  1
GN2  0  1     16  0  1
*
EREF 98 0     28  0  1
EP   97 0     99  0  1
EM   51 0     50  0  1
*
* VOLTAGE NOISE SOURCE
*
DN1  35 10    DEN
DN2  10 11    DEN
VN1  35  0    DC 2
VN2  0  11    DC 2
*
* CURRENT NOISE SOURCE
*
DN3  12 13    DIN
DN4  13 14    DIN
VN3  12  0    DC 2
VN4  0  14    DC 2
*
* CURRENT NOISE SOURCE
*
DN5  15 16    DIN
DN6  16 17    DIN
VN5  15  0    DC 2
VN6  0  17    DC 2
*
* GAIN STAGE & DOMINANT POLE AT 0.439 HZ
*
R7  18 98     1.45E7
C3  18 98     25E-9
G1  98 18     5  6  5.15E-3
V2  97 19     1.5
V3  20 51     1.5
D3  18 19     DX
D4  20 18     DX
*
* POLE/ZERO PAIR AT 1.5MHz/12.7MHz
*
R8  21 98     1E3
R9  21 22     1.25E3
C4  22 98     10E-12
G2  98 21     18 28  1E-3
*
* POLE AT 2568 MHz
*
R10 23 98     1
C5  23 98     62E-12
G3  98 23     21 28  1
*
* POLE AT 2568 MHz
*
R11 24 98     1
C6  24 98     62E-12
G4  98 24     23 28  1
*
* POLE AT 2568 MHz
*
R14 27 98     1
C8  27 98    62E-12  
G5  98 27     24 28  1
*
* COMMON-MODE GAIN NETWORK WITH ZERO AT 1 kHZ
*
R12 25 26     1E6
C7  25 26     159.155E-12
R13 26 98     1
E2  25 98      POLY(2) 1 98 2 98 0 0.28 0.28
*
*PSRR=121dB
EPSY 98 72 POLY(1) (99,50) 0 1
RPS3 72 73 1E6
CPS3 72 73 3E-9
RPS4 73 98 1
 
* OUTPUT STAGE
*
R15 28 99     100E3
R16 28 50     100E3
C9  28 50     1E-6
ISY 99 50     250E-6
R17 29 99     100
R18 29 50     100
L2  29 34     1E-9
G6  32 50     27 29  10E-3
G7  33 50     29 27  10E-3
G8  29 99     99 27  10E-3
G9  50 29     27 50  10E-3
V4  30 29     1.3
V5  29 31     3.8
F1  29  0     V4  1
F2  0  29     V5  1
D5  27 30     DX
D6  31 27     DX
D7  99 32     DX
D8  99 33     DX
D9  50 32     DY
D10 50 33     DY
*
* MODELS USED
*
.MODEL QX PNP(BF=5E5)
.MODEL DX   D(IS=1E-12)
.MODEL DY   D(IS=1E-15 BV=50)
.MODEL DZ   D(IS=1E-15 BV=7.0)
.MODEL DEN  D(IS=1E-12 RS=6.8E3 KF=1.95E-15 AF=1)
.MODEL DIN  D(IS=1E-12 RS=77.3E-6 KF=3.38E-15 AF=1)
.ENDS OP2177

