*****************
* This model was developed for Analog Devices by:
* AEI Systems, LLC
* 5777 W. Century Blvd., Suite 876
* Los Angeles, California  90045-5677
*
* The model is �2006, AEi Systems, LLC. All rights reserved. 
*
* Users may not directly or indirectly display, re-sell or 
* re-distribute this model or any derivative work therefore 
* without the prior written consent of both AEi Systems and 
* Analog Devices. This model is subject to change without 
* notice. Neither Analog Devices nor AEi Systems is responsible 
* for updating this model.
*
* For more information regarding modeling services, model 
* libraries and simulation products, please call AEi Systems 
* at (310) 216-1144, or contact AEi Systems by 
* email: info@aeng.com. Or visit AEi Systems on the web 
* at http://www.AENG.com
*$
.SUBCKT AD736 CC VIN CF NVS COM VS VOUT CAV 
* Use .OPTIONS GMIN=5E-17 for best output accuracy
R1 18 13 8K
R3 18 1 4K
R4 1 15 3K
Q1 VS 4 15 NPN
.MODEL NPN NPN
R90 6 13 3K
GB3 COM CAV VALUE={I(V4)*I(V4)}
R5 10 NVS 8K
V5 CAV 10
X3 CF COM 16 VS NVS AEIOPAMP0 
R7 CF 16 8K
R8 CC 19 8K
*R11 19 0 1G
R10 16 VOUT 0.2
GB2 VIN 0 VALUE={1P + 50P*V(VIN)}
Q7 VS 4 6 NPN
V4 13 COM
X1 1 COM 4 VS NVS AEIOPAMP1 
GB4 19 0 VALUE={1P + 15P*V(CC)}
GB1 CF COM VALUE={SQRT(I(V5))}
EB5 18 0 VALUE={IF(ABS(V(VIN)) >=ABS(V(CC)), V(VIN) , V(CC))}
.ENDS
*$
.SUBCKT AEIOPAMP0 2    3  6   7   4
RP 4 7 10K
IB 3 90 1.0000N
VIB 90 4
IO 3 2 2.5000N
RIP 3 4 1G
CIP 3 4 1.4PF
FIBN 2 4 VIB 1
RIN 2 4 1G
CIN 2 4 1.4PF
VOFST 2 10 10.0000N
RID 10 3 1G
EA 11 4 10 3 1
R1 11 12 5K
R2 12 13 50K
C1 12 4 130.00F
GA 4 14 4 13 270.00 
C2 13 14 27.000F
RO 14 4A 75
EBAL 4A 4 2A 4 1
RBAL1 7 2A 1MEG
RBAL2 2A 4 1MEG
L 14 6 300.00N
RL 14 6 1000
CL 6 4 3PF
D1 6 70 DN
VSAT 70 7 -2.0600 
D2 40 6 DN
VSAT2 40 4 2.0600 
.MODEL DN D
.ENDS
*$
.SUBCKT AEIOPAMP1 2    3  6   7   4
RP 4 7 10K
IB 3 90 5.0000N
VIB 90 4
IO 3 2 500.00P
RIP 3 4 1G
CIP 3 4 1.4PF
FIBN 2 4 VIB 1
RIN 2 4 1G
CIN 2 4 1.4PF
VOFST 2 10 10.0000N
RID 10 3 1G
EA 11 4 10 3 1
R1 11 12 5K
R2 12 13 50K
C1 12 4 65.000F
GA 4 14 4 13 135.00 
C2 13 14 13.500F
RO 14 4A 75
EBAL 4A 4 2A 4 1
RBAL1 7 2A 1MEG
RBAL2 2A 4 1MEG
L 14 6 150.00N
RL 14 6 1000
CL 6 4 3PF
D1 6 70 DN
VSAT 70 7 -1.0000 
D2 40 6 DN
VSAT2 40 4 1.0000 
.MODEL DN D
.ENDS
*$
