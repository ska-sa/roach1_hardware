* OP292 SPICE Macro-model               Rev. B, 3/95
*                                       ARG / ADSC
*
* Copyright 1993 by Analog Devices
*
* Refer to "README.DOC" file for License Statement. Use of
* this model indicates your acceptance of the terms and pro-
* visions in the License Statement.
*
* Node assignments
*                non-inverting input
*                |  inverting input
*                |  |  positive supply
*                |  |  |  negative supply
*                |  |  |  |  output
*                |  |  |  |  |
.SUBCKT OP292    2  1  99 50 34
*
* INPUT STAGE AND POLE AT 40MHZ
*
I1   99   4    50E-6
IOS  2    1    10E-9
EOS  2    3    POLY(1) (21,30) 1.5E-3 75
CIN  1    2    3E-12
Q1   5    1    7    QP
Q2   6    3    8    QP
R3   5    50   2E3
R4   6    50   2E3
R5   4    7    966
R6   4    8    966
C1   5    6    .995E-12
*
* GAIN STAGE
*
EREF 98   0    (30,0) 1
G1   98   9    (5,6) 500E-6
R7   9    98   210.819E3
D1   9    10   DX
D2   11   9    DX
V1   99   10   .6
V2   11   50   .6
*
* ZERO/POLE AT 6MHZ/12MHZ
*
E1   12   98   (9,30) 2
R8   12   13   1
R9   13   98   1
C3   12   13   26.526E-9
*
* ZERO AT 15MHZ
*
E2   14   98   (13,30) 1E6
R10  14   15   1E6
R11  15   98   1
C4   14   15   10.610E-15
*
* COMMON MODE STAGE WITH ZERO AT 40KHZ
*
ECM  20   98   POLY(2) (1,30) (2,30) 0 0.5 0.5
R20  20   21   1E6
R21  21   98   1
C5   20   21   3.979E-12
*
* POLE AT 100MHZ
*
G2   98   16   (15,30) 1
R12  16   98   1
C6   16   98   1.592E-9
*
* OUTPUT STAGE
*
RS1  99   30   1E6
RS2  30   50   1E6
ISY  99   50   .44E-3
G3   31   50   POLY(1) (16,30) -1.635E-6 4E-6
R16  31   50   1E6
DCL  50   31   DZ
I2   99   32   250E-6
RCL  33   50   56
M1   32   31   50   50   MN L=9E-6 W=1000E-6 AD=15E-9 AS=15E-9
M2   34   31   50   50   MN L=9E-6 W=1000E-6 AD=15E-9 AS=15E-9
CC   31   32   14E-12
Q3   99   32   34   QNA
Q4   33   32   34   QPA
Q5   31   33   50   QNA
.MODEL QNA NPN(IS=1.19E-16 BF=253 NF=0.99 VAF=193 IKF=2.76E-3
+ ISE=2.57E-13 NE=5 BR=0.4 NR=0.988 VAR=15 IKR=1.465E-4
+ ISC=6.9E-16 NC=0.99 RB=2.0E3 IRB=7.73E-6 RBM=132.8 RE=4 RC=209
+ CJE=2.1E-13 VJE=0.573 MJE=0.364 FC=0.5 CJC=1.64E-13 VJC=0.534 MJC=0.5
+ CJS=1.37E-12 VJS=0.59 MJS=0.5 TF=0.43E-9 PTF=30)
.MODEL QPA PNP(IS=5.21E-17 BF=131 NF=0.99 VAF=62 IKF=8.35E-4
+ ISE=1.09E-14 NE=2.61 BR=0.5 NR=0.984 VAR=15 IKR=3.96E-5
+ ISC=7.58E-16 NC=0.985 RB=1.52E3 IRB=1.67E-5 RBM=368.5 RE=6.31 RC=354.4
+ CJE=1.1E-13 VJE=0.745 MJE=0.33 FC=0.5 CJC=2.37E-13 VJC=0.762 MJC=0.4
+ CJS=7.11E-13 VJS=0.45 MJS=0.412 TF=1.0E-9 PTF=30) 
.MODEL MN NMOS(LEVEL=3 VTO=1.3 RS=0.3 RD=0.3 
+ TOX=8.5E-8 LD=1.48E-6 WD=1E-6 NSUB=1.53E16 UO=650 DELTA=10 VMAX=2E5
+ XJ=1.75E-6 KAPPA=0.8 ETA=0.066 THETA=0.01 TPG=1 CJ=2.9E-4 PB=0.837
+ MJ=0.407 CJSW=0.5E-9 MJSW=0.33)
.MODEL QP PNP(BF=61.5)
.MODEL DX D
.MODEL DZ D(BV=3.6)
.ENDS
