* AD9624 SPICE MACRO MODEL                  3/94, REV. B
*   CLD
*
* Revision History:
*     Changed parameter VJ=-1 to VJ=0.01 in diode model. 
*
* Copyright 1992 by Analog Devices, Inc.
*
* Refer to "README.DOC" file for License Statement.  Use of this model
* indicates your acceptance with the terms and provisions in the License Statement.
*
*
* NODE ASSIGNMENTS
*              POSITIVE INPUT
*              |    NEGATIVE INPUT
*              |    |    POSITIVE SUPPLY
*              |    |    |
*              |    |    |   NEGATIVE SUPPLY
*              |    |    |   |   OUTPUT
*              |    |    |   |   |
.SUBCKT AD9624 VINP VINN 100 110 VOUT 
*
C1   5    VOUT 4E-12
C2 VOUT 6 4E-12
F1 100 5 V1 1
F2 6 110 V2 1
G1 100 9 POLY(1) (5,0) 0.392 -0.13
G2 10 110 POLY(1) (6,0) 0.392 0.13
GM1 5 7 POLY(1) (1,3) 0.005     0.025
GM2 8 6 POLY(1) (2,4) 0.005 -0.025
D1 9 100 D
D2 110 10 D
V1 100 8 0
V2 7 110 0
V3 6A 0 DC -2.4
D3 6A 6 D1
V4 5A 0 DC 2.4
D4 5 5A D1
V5 5B 0 DC 3.5
D5 5B 5 D1
V6 6B 0 DC -3.5
D6 6 6B D1
I1 100 1 .7E-3
I2 2 110 1.1E-3
I3 100 3 .7E-3
I4 4 110 1.1E-3
Q1 110 VINP 1 100 PA
Q2 100 VINP 2 110 NA
Q3 100 VINN 4 110 NA
Q4 110 VINN 3 100 PA
Q5 9 9 13 110 NB 1.2
Q6 10 10 13 100 PB
Q7 100 9 11 110 NB 2.4  
Q8 110 10 12 100 PB 2  
R1 100 5 300
R2 6 110 300
R3 5 0 450
R4 6 0 450
R5 11 VOUT 7
R6 VOUT 12 7
***
.MODEL NA NPN
 + IS   = 1.6E-16  BF   = 305 VAF  = 74
 + IKF  = 2.2E-02  ISE  = 2E-17  NE   = 1.2  BR   = 36
 + VAR  = 1.7  IKR  = 3.0E-02  ISC  = 1.5E-19 
 + NC   = 1.7  RB   = 90  IRB  = 0  RBM  = 20
 + RE   = 0.9  RC   = 52  CJE  = 1.2E-13  VJE  =0.8 
 + MJE  = 0.5  TF   = 2.8E-11  XTF  = 5.0  VTF  = 2.7 
 + ITF  = 2.6E-02  PTF  = 0.0  CJC  = 1.7E-13  VJC  = 0.6
 + MJC  = 0.34  XCJC = 0.138  TR   = 7.1E-11  CJS  = 3.9E-13 
 + VJS  = 0.5  MJS  = 0.32  XTB  = 1.1  EG   = 1.18 
 + XTI  = 2.0  FC   = 0.82 
.MODEL NB NPN
 + IS   = 6.4E-16  BF   = 305  VAF  = 74 
 + IKF  = 8.7E-02  ISE  = 8E-17  NE   = 1.2  BR   = 40 
 + VAR  = 1.7  IKR  = 0.12  ISC  = 4.6E-19 
 + NC   = 1.7  RB   = 23 IRB  = 0  RBM  = 5.0 
 + RE   = 0.227  RC   = 9.5  CJE  = 4.8E-13  VJE  = 0.8 
 + MJE  = 0.5  TF   = 2.7E-11  XTF  = 5.1  VTF  = 2.7 
 + ITF  = 0.11  PTF  = 0.0  CJC  = 5.0E-13  VJC  = 0.60
 + MJC  = 0.34  XCJC = 0.19  TR   = 7.1E-11  CJS  = 6.9E-13 
 + VJS  = 0.5  MJS  = 0.32  XTB  = 1.1  EG   = 1.18 
 + XTI  = 2.0  FC   = 0.82 
.MODEL PA PNP
 + IS   = 6.3E-17  BF   = 69  VAF  = 25 
 + IKF  = 9.1E-03  ISE  = 3.2E-16  NE   = 1.4  BR   = 16 
 + VAR  = 1.8  IKR  = 6.7E-02  ISC  = 1.9E-18 
 + NC   = 1.6  RB   = 57  IRB  = 0  RBM  = 15 
 + RE   = 1.3  RC   = 51  CJE  = 8.0E-14  VJE  = 0.82 
 + MJE  = 0.49  TF   = 2.6E-11  XTF  = 9.0  VTF  = 2.7 
 + ITF  = 2.7E-02  PTF  = 0.0  CJC  = 2.4E-13  VJC  = 0.53 
 + MJC  = 0.19  XCJC = 0.13  TR   = 6.5E-11  CJS  = 6.9E-13 
 + VJS  = 0.60  MJS  = 0.35  XTB  = 2.5 EG   = 1.18 
 + XTI  = 2.0  FC   = 0.90 
.MODEL PB PNP
 + IS   = 3.8E-16  BF   = 69  VAF  = 25 
 + IKF  = 5.5E-02  ISE  = 1.9E-15  NE   = 1.4  BR   = 19 
 + VAR  = 1.8  IKR  = 0.4  ISC  = 1.1E-17 
 + NC   = 1.6  RB   = 9.5  IRB  = 0  RBM  = 2.5 
 + RE   = 0.21  RC   = 15  CJE  = 4.8E-13  VJE  = 0.82 
 + MJE  = 0.49E-01  TF   = 2.4E-11  XTF  = 9.0  VTF  = 2.7 
 + ITF  = 0.16  PTF  = 0.0  CJC  = 9.5E-13  VJC  = 0.53 
 + MJC  = 0.19  XCJC = 0.19  TR   = 6.5E-11  CJS  = 1.5E-12 
 + VJS  = 0.6  MJS  = 0.35  XTB  = 2.5  EG   = 1.18 
 + XTI  = 2.0  FC   = 0.9 
.MODEL D D (CJO=30E-12 VJ=0.01 M=2 )  
.MODEL D1 D (IS=1E-14 )  
.ENDS
*
* TEST CIRCUIT
*
*VIN VINPA 0 DC 0 AC 1 PULSE(-.3125 .3125  5.000n 2.000n 2.000n 30.000n 65.000n ) 
*VIN VINPA 0 DC 0 AC 1 SIN (0 .125 20MEG 0 0 0)
*VCC 100 0 DC 5 AC 0
*VEE 110 0 DC -5 AC 0
*RT VINPA VINP 25
*RL VOUT 0 100
*RF VOUT VINN 430
*RN VINN 0 62
*
*X1 VINP VINN 100 110 VOUT AD9624
*
*.END
