* AD8502 SPICE Macro-model
* Typical Values
* 14 May 2007, Version 1.0
* HH ADSJ
*
* Copyright 2007 by Analog Devices
*
* Refer to "README.DOC" file for License Statement.  Use of this
* model indicates your acceptance of the terms and provisions in
* the License Statement.
*
* Node Assignments
*                       noninverting input
*                       |   inverting input
*                       |   |    positive supply
*                       |   |    |   negative supply
*                       |   |    |   |   output
*                       |   |    |   |   |
*                       |   |    |   |   |
.SUBCKT AD8502          1   2   99  50  45
*
* INPUT STAGE
*
MI1  14  7  8  8 PIX 
MI2  16  2  8  8 PIX
MI3  17  7 10 10 NIX
MI4  18  2 10 10 NIX
RD1 14 50 1.33E+06
RD2 16 50 1.33E+06
RD3 99 17 1.33E+06
RD4 99 18 1.33E+06
C1  14 16 4.53E-12
C2  17 18 4.53E-12
I1  99  8 3.00E-07
I2  10 50 3.00E-07
V1  99  9 0.220E+00
V2  13 50 0.220E+00
D1   8  9 DX
D2  13 10 DX
EOS  7  1 POLY(4) (22,98) (73,98) (81,98) (70,98) 5.00E-04 1 1 1 1
IOS  1  2 2.50E-13
*
*CMRR=100dB, POLE AT 12 Hz
*
E1  21 98 POLY(2) (1,98) (2,98) 0 8.33E-03 8.33E-03
R10 21 22 1.33E+04
R20 22 98 7.96E-01
C10 21 22 1.00E-06
*
* PSRR=80dB, POLE AT 5 Hz
*
EPSY 72 98 POLY(1) (99,50) -125.00  25.00
CPS3 72 73 1.00E-06
RPS3 72 73 3.98E+04
RPS4 73 98 1.59E-01
*
* VOLTAGE NOISE REFERENCE OF 190nV/rt(Hz)
*
VN1 80 98 0
RN1 80 98 16.45E-3
HN  81 98 VN1 1.74E+02
RN2 81 98 1
*
* FLICKER NOISE CORNER = 7 Hz
*
D5  69 98 DNOISE
VSN 69 98 DC 0.6551
H1  70 98 POLY(1) VSN 1.00E-03 1.00E+00
RN  70 98 1
*
* INTERNAL VOLTAGE REFERENCE
*
EREF 98  0 POLY(2) (99,0) (50,0) 0 0.5 0.5
GSY  99 50 POLY(1) (99,50) +1E-10 1.95E-08
EVP  97 98 POLY(1) (99,50) 0 0.5
EVN  51 98 POLY(1) (50,99) 0 0.5
*
* GAIN STAGE
*
G1 98 30 POLY(2) (14,16) (17,18) 0 2.54E-07 2.54E-07
R1 30 98 1.00E+06
RZ 30 31 1.00E-03
CF 45 31 5.08E-11

V3 32 30  0.495E+00
V4 30 33  0.281E+00
D3 32 97 DX
D4 51 33 DX
*
* OUTPUT STAGE
*
MO5  45 46 99 99 POX  
MO6  45 47 50 50 NOX 
EG1 99 46 POLY(1) (98,30)  6.024E-01 1 ;  PMOS
EG2 47 50 POLY(1) (30,98)  6.012E-01 1 ;  NMOS 
*
* MODELS
*
.MODEL POX PMOS (LEVEL=2,KP=5.00E-05,VTO=-0.6,LAMBDA=0.03,RD=0, L=1.0E-6, W=1.10E-03,RD=0)
.MODEL NOX NMOS (LEVEL=2,KP=5.00E-05,VTO=+0.6,LAMBDA=0.03,RD=0, L=1.0E-6, W=4.63E-03, RD=0)
.MODEL PIX PMOS (LEVEL=2,KP=5.00E-05,VTO=-0.5,LAMBDA=0.03, L=1E-6, W=9.31E-07)
.MODEL NIX NMOS (LEVEL=2,KP=5.50E-05,VTO=0.5,LAMBDA=0.03, L=1E-6, W=9.31E-07)
.MODEL DX D(IS=1E-14,RS=5)
.MODEL DNOISE D(IS=1E-14,RS=0,KF=8.53E-11)
*
*
.ENDS AD8502
*
*$
