* OP186 SPICE Macro-model Typical Values
* 2/98, Ver. 1
* TAM / ADSC
*
* Copyright 1998 by Analog Devices
*
* Refer to "README.DOC" file for License Statement.  Use of this
* model indicates your acceptance of the terms and provisions in
* the License Statement.
*
* Node Assignments
*			noninverting input
*			|	inverting input
*			|	|	 positive supply
*			|	|	 |	 negative supply
*			|	|	 |	 |	 output
*			|	|	 |	 |	 |
*			|	|	 |	 |	 |
.SUBCKT OP186		1	2	99	50	45
*
* INPUT STAGE
*
Q1   4  1 3 PIX
Q2   6  7 5 PIX
RC1  4 50 100E3
RC2  6 50 100E3
RE1  3  8 6.452E3
RE2  5  8 6.452E3
C1   4  6 50E-15
I1  99  8 1E-6
EOS  7  2 POLY(2) (12,98) (73,98) 800E-6 1 1
IOS  1  2 50E-12
V1  99  9 0.9
V2  99 10 0.9
D1   3  9 DX
D2   5 10 DX
*
* CMRR 90dB, ZERO AT 1kHz
*
ECM1 11 98 POLY(2) (1,98) (2,98) 0 .5 .5
RCM1 11 12 1.59E6
CCM1 11 12 100E-12
RCM2 12 98 50
*
* PSRR=100dB, ZERO AT 200Hz
*
RPS1 70  0 1E6
RPS2 71  0 1E6
CPS1 99 70 1E-5
CPS2 50 71 1E-5
EPSY 98 72 POLY(2) (70,0) (0,71) 0 1 1
RPS3 72 73 1.59E6
CPS3 72 73 500E-12
RPS4 73 98 15.9
*
* INTERNAL VOLTAGE REFERENCE
*
* RSY1 99 91 10E6
* RSY2 50 90 10E6
* VSN1 91 90 DC 0
* EREF 98  0 (90,0) 1
EREF 98  0 POLY(2) (99,0) (50,0) 0 .5 .5
GSY  99 50 POLY(1) (99,50) 2E-6 .1E-6
*
* POLE AT 600kHz; ZERO AT 900kHz
*
G1 98 20 (4,6) 11.3E-6
R1 20 98 88.46E3
R2 20 21 176.8E3
C2 21 98 1E-12
*
* GAIN STAGE
*
G4  98 30 (20,98) 19.54E-6
R7  30 98 111.6E6
CF  45 30 32E-12
D3  30 31 DX
D4  32 30 DX
V3  99 31 0.6
V4  32 50 0.6
*
* OUTPUT STAGE
*
M1  45 46 99 99 POX L=2u W=100u
M2  45 47 50 50 NOX L=2u W=98u
EG1 99 46 POLY(1) (98,30) 0.82 1
EG2 47 50 POLY(1) (30,98) 0.79 1
*
* MODELS
*
.MODEL POX PMOS (LEVEL=2, KP=10E-6, VTO=-0.75, LAMBDA=0.01)
.MODEL NOX NMOS (LEVEL=2, KP=17E-6, VTO=0.75,  LAMBDA=0.01)
.MODEL PIX PNP (BF=185,KF=1.6E-12,AF=1)
* .MODEL PIX2 PNP (BF=200,IS=1E-16)
.MODEL DX D(IS=1E-14)
.ENDS OP186