* OP250/OP450 SPICE Macro-Model Typcial Values
* 10/97, Ver. 1
* TAM / ADSC
*
* Node assignments
*		noninverting input
*		|	inverting input
*		|	|	positive supply
*		|	|	|	negative supply
*		|	|	|	|	output
*		|	|	|	|	|
*		|	|	|	|	|
.SUBCKT OP250	1	2	99	50	45
*
* INPUT STAGE
*
M1  4  3  6 6 MNIN L=2u W=66u
M2  5  2  6 6 MNIN L=2u W=66u
M3  7  3  9 9 MPIN L=2u W=66u
M4  8  2  9 9 MPIN L=2u W=66u
RD1   99  4 5E3
RD2   99  5 5E3
RD3    7 50 5E3
RD4    8 50 5E3
VCM1  10 50 -.3
VCM2  99 11 -.3
D1    10  6 DX
D2     9 11 DX
EOS    3  1 POLY(3) (61,98) (73,98) (81,0) 3E-3 1 1 1
IOS    1  2 .25E-12
IBIAS1  6 50 700E-6
IBIAS2 99  9 700E-6
*
* CMRR=60 dB, ZERO AT 20kHz
*
ECM1 60 98 POLY(2) (1,98) (2,98) 0 .5 .5
RCM1 60 61 159.2E3
RCM2 61 98 159
CCM1 60 61 50E-12
*
* PSRR=90dB, ZERO AT 200Hz
*
RPS1 70  0 1E6
RPS2 71  0 1E6
CPS1 99 70 1E-5
CPS2 50 71 1E-5
EPSY 98 72 POLY(2) (70,0) (0,71) 0 1 1
RPS3 72 73 1.59E6
CPS3 72 73 500E-12
RPS4 73 98 50
*
* INTERNAL VOLTAGE REFERENCE
*
RSY1 99 91 100E3
RSY2 50 90 100E3
VSN1 91 90 DC 0
EREF 98  0 (90,0) 1
GSY  99 50 POLY(1) (99,50) -1.81E-3 1.5E-5
*
* VOLTAGE NOISE REFERENCE OF 30nV/rt(Hz)
*
VN1 80 0 0
RN1 80 0 16.45E-3
HN  81 0 VN1 30
RN2 81 0 1
*
* POLE AT 1.25MHz
*
G2 98 20 POLY(2) (4,5) (7,8) 0 5E-5 5E-5
R2 20 98 10E3
C2 20 98 12.7E-12
*
* GAIN STAGE
*
G1 98 30 (20,98) 3.5E-4
R1 30 98 6.25E6
CF 30 45 135E-12
D4 31 99 DX
D5 50 32 DX
V1 31 30 0.7
V2 30 32 0.7
*
* OUTPUT STAGE
*
M5  45 41 99 99 MPOUT L=2u W=6660u
M6  45 42 50 50 MNOUT L=2u W=6660u
EO1 99 41 POLY(1) (98,30) .9232 1
EO2 42 50 POLY(1) (30,98) .8914 1
*
* MODELS
*
.MODEL MNIN  NMOS(LEVEL=2,VTO=0.75,KP=20E-6,CGSO=0,KF=2.5E-31,AF=1)
.MODEL MPIN  PMOS(LEVEL=2,VTO=-0.75,KP=20E-6,CGSO=0,KF=2.5E-31,AF=1)
.MODEL MNOUT NMOS(LEVEL=2,VTO=0.75,KP=30E-6,LAMBDA=0.04,CGSO=0)
.MODEL MPOUT PMOS(LEVEL=2,VTO=-0.75,KP=20E-6,LAMBDA=0.04,CGSO=0)
.MODEL DX D(IS=1E-16)
.ENDS OP250