* REF43 SPICE MACROMODEL                     4/96, Rev. A
*                                            (RN)  
*
* 
*
* Refer to "README.DOC" file for License Statement.  Use of this
* model indicates your acceptance with the terms and provisions in
* the License Statement.
*
*  NODE NUMBERS
*               VIN
*               |  GND
*               |  |  TRIM
*               |  |  |  VOUT
*               |  |  |  |
.SUBCKT REF43   2  4  5  6
*
* 1.23V REFERENCE
*
I1     4  10   1.22998E-3
R1     10  4   1E3  TC=6E-6
EN     10  9   41 0  1
G1     4   9   2  4  983.9E-12
F1     4   9   VS  17.0565E-6
*
* NOISE GENERATOR
*
VN1    40  0   DC  2
DN1    40  41  DEN
DN2    41  42  DEN
VN2    0   42  DC  2
*
* INTERNAL OP AMP
*
G2     4  11   9  19  1E-3
R2     4  11   300E6
C1     4  11   5E-10
D1     11 12   DX
V1     2  12   1.5
*
* SECONDARY POLE
*
G3     4  13   11 4  1E-6
R3     4  13   1E6
C2     4  13   1.5E-13
*
* OUTPUT STAGE
*
ISY    2   4   0.246E-3
FSY    2   4   V1  -1 
G4     4  14   13  4  25E-6
R4     4  14   40E3
R7     17 19   13.6E3
R8     19  4   13.1716E3
R9     19  5   196E3
R10    5   4   1E12
Q1     16 14   17   QN
VS     18 17   DC 0
L1     18  6   1E-9
*
* OUTPUT CURRENT LIMIT
*
Q2     15  2   16  QN
R6     2  16   14
R5     2  15   18E3
C3     2  15   1E-6
G5     14  4   2  15  1
*

.MODEL  QN  NPN(IS=1E-15  BF=1000)
.MODEL  DX  D(IS=1E-15)
.MODEL  DEN D(IS=1E-12 RS=1.3796e6 AF=1 KF=1.998751E-17)
.ENDS
