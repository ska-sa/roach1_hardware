* OP279 SPICE Macro-model               Rev. A, 7/94
*                                       ARG / PMI
*
* Copyright 1994 by Analog Devices
*
* Refer to "README.DOC" file for License Statement. Use of
* this model indicates your acceptance of the terms and pro-
* visions in the License Statement.
*
* Node assignments
*                non-inverting input
*                |  inverting input
*                |  |  positive supply
*                |  |  |  negative supply
*                |  |  |  |  output
*                |  |  |  |  |
.SUBCKT OP279    3  2  99 50 45
*
* INPUT STAGE AND POLE AT 6MHZ
*
I1   1    50   60.2E-6
Q1   5    2    7    QN
Q2   6    4    8    QN
D1   4    2    DX
D2   2    4    DX
R1   1    7    1.628E3
R2   1    8    1.628E3
R3   5    99   2.487E3
R4   6    99   2.487E3
C1   5    6    5.333E-12
EOS  4    3    POLY(1) (16,39) 0.25E-3 50.118
IOS  2    3    5E-9
GB1  2    98   (24,98) 100E-9
GB2  4    98   (24,98) 100E-9
CIN  2    3    1E-12
*
* GAIN STAGE AND DOMINANT POLE AT 16HZ
*
EREF 98   0    (39,0) 1
G1   98   9    (5,6) 402.124E-6
R7   9    98   497.359E6
C2   9    98   20E-12
V1   99   10   0.58
V2   11   50   0.47
D5   9    10   DX
D6   11   9    DX
*
* COMMON MODE STAGE WITH ZERO AT 10KHZ
*
ECM  15   98   POLY(2) (3,39) (2,39) 0 0.5 0.5
R9   15   16   1E6
R10  16   98   10
C3   15   16   15.915E-12
*
* ZERO AT 1.5MHZ
*
E1   14   98   (9,39) 1E6
R5   14   18   1E6
R6   18   98   1
C4   14   18   106.103E-15
*
* BIAS CURRENT-VS-COMMON MODE VOLTAGE
*
EP   97   0    (99,0) 1
EN   51   0    (50,0) 1
V3   20   21   1.6
V4   22   23   2.8
R12  97   20   530
R13  23   51   1E3
D13  15   21   DX
D14  22   15   DX
FIB  98   24   POLY(2) V3 V4 0 -1 1
RIB  24   98   10E3
E3   97   25   POLY(1) (99,39) -1.63 1
E4   26   51   POLY(1) (39,50) -2.73 1
D15  24   25   DX
D16  26   24   DX
*
* POLE AT 6MHZ
*
G6   98   40   (18,39) 1E-6
R20  40   98   1E6
C10  40   98   26.526E-15
*
* OUTPUT STAGE
*
RS1  99   39   6.0345E3
RS2  39   50   6.0345E3
RO1  99   45   40
RO2  45   50   40
G7   45   99   (99,40) 25E-3
G8   50   45   (40,50) 25E-3
G9   98   60   (45,40) 25E-3
D9   60   61   DX
D10  62   60   DX
V7   61   98   DC 0
V8   98   62   DC 0
FSY  99   50   POLY(2) V7 V8 1.711E-3  1  1
D11  41   45   DZ
D12  45   42   DZ
V5   40   41   1.54
V6   42   40   1.54
.MODEL DX D()
.MODEL DZ D(IS=1E-6)
.MODEL QN NPN(BF=300)
.ENDS
