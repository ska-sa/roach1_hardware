* AD8004a SPICE Macro-model                  12/96, revA
*                                           SMR/ADI
*
* Copyright 1996 by Analog Devices, Inc.
*
* Refer to "README.DOC" file for License Statement.  Use of this model
* indicates your acceptance with the terms and provisions in the License Statement.
*
* This model was written with the specs as they apply to running from a
* dual supply, +/-5v. This means that the model will give a slew rate of
* 3000v/us, whether or not the model is run from +/-5v, or single supply
* of 5v. The user should keep in mind that the actual slew rate is much 
* slower in the real device when running from single supply 5v. Refer to
* the data sheet for the actual specs. 
*
* Node assignments
*                non-inverting input
*                | inverting input
*                | | positive supply
*                | | |  negative supply
*                | | |  |  output
*                | | |  |  |
.SUBCKT AD8004a  1 2 99 50 24   
*
* INPUT STAGE
*
r1   99 8 1
r2   10 50 1
i1   99 5 100e-6
i2   4 50 100e-6
q1   50 3 5  qp1
q2   99 3 4  qn1
q3   8 6 2  qn2
q4   10 7 2 qp2
r3   5 6 1
r4   4 7 1
r3a  99 6 40k
r4a  50 7 40k
*
* input error sources
* 
ib1  99  2     90e-6
ib2  99  3     110e-6
vos  3   1     3.5e-3
cs1  99  2     0.75e-12
cs2  50  2     0.75e-12
cs3  99  3     0.75e-12
cs4  50  3     0.75e-12
*
* first gain stage and dominant pole
*
r5   12 99     280k
r6   12 50     280k
c3   12 99     1e-12
c4   12 50     1e-12
g1   99 12     99 8 1
g2   12 50     10 50 1 
gsl1 99 12     poly(1) 99 8 0 0 300
gsl2 12 50     poly(1) 10 50 0 0 300
v3   99 13     1.6
v4   14 50     1.6
d3   12 13     dx
d4   14 12     dx
*
* secondary pole
*
r7  15 99    1k
r8  15 50    1k
c5  15 99    0.9pf
c6  15 50    0.9pf
g3  99 15    12 18 1e-3
g4  15 50    18 12 1e-3
*
* buffer stage
*
g13 98 17 15 98 1e-4    
rbuf 17 98 10k
*
* reference stage
*
r13 18 99 1e5 
r14 18 50 1e5
eref 98 0 18 0 1 
rref 98 0 1e6
*
* current mirroring on supplies
*
fo1 98 300 vcd 1
vi1 311 98 0
vi2 98 312 0
dm1 300 311 dx
dm2 312 300 dx
fsy 99 50 poly(2) vi1 vi2 0 1 1
iq 99 50 10.9e-3
*
* output stage
*
r15 23 99   2
r16 23 50   2
vcd 23 25   0
l1  25 24   1.5e-12
rl  24 98   1e6
g11 99 23   17 99  0.5
g12 23 50   50 17  0.5
v5  19 23   0.59
v6  23 20   0.59
d5  19 17   dx
d6  17 20   dx
*
* models
*
.model qn1 npn(bf=1e3 is=1e-15)
.model qp1 pnp(bf=1e3 is=1e-15)
.model qn2 npn(bf=1e3 is=1e-15)
.model qp2 pnp(bf=1e3 is=1e-15)
.model dx   d(is=1e-15)
.ends ad8004a
