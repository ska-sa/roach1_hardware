* AD848 SPICE Macro-model                   3/94, Rev. B
*                                           JCB / PMI
*
* Revision History:
*     Changed Negative Zero stage to remove the
*     negative capacitor value. 
*
* Copyright 1990 by Analog Devices
*
* Refer to "README.DOC" file for License Statement.
* Use of this model indicates your acceptance with the
* terms and provisions in the License Statement.
*
* Node assignments
*               non-inverting input
*               | inverting input
*               | | positive supply
*               | | |  negative supply
*               | | |  |  output
*               | | |  |  |
*               | | |  |  |
.SUBCKT AD848   1 2 99 50 30
*
* INPUT STAGE & POLE AT 400 MHZ
*
R1   2  3     5E11
R2   1  3     5E11
R3   5 99     62.5
R4   6 99     62.5
CIN  1  2     1.5E-12
C2   5  6     3.184E-12
I1   4  50    4.0E-3
IOS  1  2     25E-9
EOS  9  1     POLY(1)  20 23  0.5E-3  1
Q1   5  2 10  QX
Q2   6  9 11  QX
R5   10 4     49.6
R6   11 4     49.6
*
EREF 98 0     23  0  1
*
* GAIN STAGE & DOMINANT POLE AT 10 KHZ
*
R7  12 98     1.25E6
C3  12 98     12.74E-12
G1  98 12     5  6  16.0E-3
V2  99 13     1.7
V3  14 50     1.7
D3  12 13     DX
D4  14 12     DX
*
* NEGATIVE ZERO AT 160 MHZ
*
R8  15 16     1E6
R9  16 98     1
FX1 15 16     VX1  -1
E1  15 98     12 23  1E6
VX1 80  0     0
EX1 81  0     15  16  1
C4  80 81     0.995E-15
*
* POLE AT 400 MHZ
*
R10 17 98     1E6
C5  17 98     398E-18
G2  98 17     16 23  1E-6
*
* POLE AT 400 MHZ
*
R11 18 98     1E6
C6  18 98     398E-18
G3  98 18     17 23  1E-6
*
* COMMON-MODE GAIN NETWORK WITH ZERO AT 100 kHZ
*
R12 19 20     1E6
C7  19 20     1.59E-12
R13 20 98     1
E2  19 98     3  23  5.62
*
* POLE AT 400 MHZ
*
R14 21 98     1E6
C8  21 98     398E-18
G4  98 21     18 23  1E-6
*
* OUTPUT STAGE
*
RF  25 22     500
CF  22 12     12.5E-12
R16 23 99     25E3
R17 23 50     25E3
ISY 99 50     0.5E-3
R18 25 99     90
R19 25 50     90
L2  25 30     3E-8
G5  28 50     21 25  11.11E-3
G6  29 50     25 21  11.11E-3
G7  25 99     99 21  11.11E-3
G8  50 25     21 50  11.11E-3
V4  26 25     0.8
V5  25 27     0.8
D5  21 26     DX
D6  27 21     DX
D7  99 28     DX
D8  99 29     DX
D9  50 28     DY
D10 50 29     DY
*
* MODELS USED
*
.MODEL QX NPN(BF=606.1)
.MODEL DX   D(IS=1E-15)
.MODEL DY   D(IS=1E-15 BV=50)
.ENDS
