* AMP01 SPICE Macro-model                 2/90, Rev. A
*                                          DFB / PMI
*
* Copyright 1990 by Analog Devices, Inc.
*
* Refer to "README.DOC" file for License Statement.  Use of this model
* indicates your acceptance with the terms and provisions in the License Statement.
*
* Node assignments
*
*              rg(pin1)
*              |   rg(pin2)
*              |   |   inverting input
*              |   |   | sense
*              |   |   | |   reference
*              |   |   | |   |   output
*              |   |   | |   |   |                              
.SUBCKT AMP01  207 206 2 210 209 32 211 50 99 212 214 216 3
*                                   |   |  |  |   |   |   |
*        output stage negative supply   |  |  |   |   |   |
*                 device negative supply   |  |   |   |   |
*                     device positive supply  |   |   |   |
*                  output stage positive supply   |   |   |
*                                                rs   |   |
*                                                    rs   |
*                                       non-inverting input
*input protection network
*
R201 3 204 250
R202 2 205 250
D202 206 204 DX
D203 207 205 DX
*
*input stage and resistive load
*
Q201 6 204 206 NX
Q202 5 205 207 NX
R3 99 6 30K
R4 99 5 30K
*
*common mode rejection term
*
R207 99 207 8E12
R208 50 207 8E12
*
*input offset current and input offset voltage
*
I202 99 204 150E-9
I203 3 50 149.5E-9
*
*output offset voltage
*
I201 99 201 40E-9
*
*feedback V-I converter
*
C2 201 202 120E-12
*c2 provides the second pole before the
*input stage to prevent spurious slew limiting
R203 209 201 47.5K
R204 201 203 2.5K
R205 202 203 2.5K
R206 210 202 47.5K
V203 203 50 0.57
E201 213 50 201 214 100K
Q203 206 213 214 NX
I204 214 50 100E-6
E202 215 50 202 216 100K
Q204 207 215 216 NX
I205 216 50 100E-6
D204 208 207 DX
D205 208 206 DX
V201 208 50 4
*
* output amplifier
*
R5 9 99 400E6
R6 9 50 400E6
C3 9 99 55E-12
C4 9 50 55E-12
G1 99 9 POLY(1) 5 6 1.7M 100E-6
G2 9 50 POLY(1) 6 5 1.7M 100E-6
V2 99 8 2.5
V3 10 50 2.5
D1 9 8 DX
D2 10 9 DX
D5 9 28 DX
D6 29 9 DX
R26 26 212 111E3
R27 26 211 111E3
R28 32 212 90
R29 32 211 90
G17 30 211 9 32 11.111E-3
G18 31 211 32 9 11.111E-3
G19 32 212 212 9 11.111E-3
G20 211 32 9 211 11.111E-3
V6 28 32 3
V7 32 29 3
D7 212 30 DX
D8 212 31 DX
D9 211 30 DY
D10 211 31 DY
I1 212 211 600E-6
*
* non-linear models
*
.MODEL DX D (IS=1E-15)
.MODEL DY D (IS=1E-15 BV=50)
.MODEL NX NPN (IS=1E-14 BF=1E5 RE=50)
.ENDS
