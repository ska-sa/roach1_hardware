* MLT04  SPICE Macro-model              Rev. A, 12/93
*                                       JCB / ADI
*
* Copyright 1993 by Analog Devices
*
* Refer to "README.DOC" file for License Statement.  Use of
* this model indicates your acceptance of the terms and pro-
* visions in the License Statement.
*
* Node assignments
*                X-input
*                |  Y-input
*                |  |  Ground
*                |  |  |  W-output
*                |  |  |  |  Positive supply
*                |  |  |  |  |  Negative supply
*                |  |  |  |  |  |
.SUBCKT MLT04    3  4  2  1  99 50
*
* X AND Y INPUT STAGES
*
V1   3   20    10.5E-3
C1   20   2    3E-12
R1   20   2    1E6
I1   20   2    2.3E-6
V2   4   21    10.5E-3
C2   21   2    3E-12
R2   21   2    1E6
I2   21   2    2.3E-6
*
* MULTIPLIER CORE
*
G1   98  22    POLY(2)  (20,2) (21,2)  (0,0,0,0,0.4E-6)
R3   98  22    1E6
C3   98  22    1E-15
*
* INPUT STAGE
*
I3   99  28    1E-4
Q1   24   1    26   QP
Q2   25  23    27   QP
R4   50  24    11635
R5   50  25    11635
R6   26  28    11119
R7   27  28    11119
E1   23  98    POLY(1) (22,98)  -10E-3  1
*
* GAIN STAGE AND DOMINANT POLE AT 145HZ
*
EREF 98  0     POLY(2) (99,0) (50,0) 0 0.5 0.5
G2   98  29    (24,25) 8.59E-5
R8   29  98    5.82E8
C4   29  98    1.89E-12
D1   29  30    DX
D2   31  29    DX
V3   99  30    2.2
V4   31  50    2.2
*
*POLE AT 30MHZ
*
G3   98  32    (29,98) 1E-6
R9   32  98    1E6
C5   32  98    5.31E-15
*
* OUTPUT STAGE
*
R10  99   1    80
R11  1   50    80
G4   1   99    (99,32) 12.5E-3
G5   50   1    (32,50) 12.5E-3
D3   32  33    DX
D4   34  32    DX
V5   33   1    0.72
V6   1   34    0.72
G6   98  35    (1,32)  12.5E-3
D5   35  36    DX
D6   37  35    DX
V7   36  98    DC 0
V8   98  37    DC 0
F1   99  50    POLY(2) V7 V8 3.65E-3  1  1
*
* MODELS USED
*
.MODEL DX D
.MODEL QP PNP(BF=143)
.ENDS