* AD840J SPICE Macro-model                 1/91, Rev. A   
*                                           AAG / PMI
*
* This version of the AD-840 model simulates the worst case 
* parameters of the 'J' grade.  The worst case parameters
* used correspond to those in the data sheet.
*
* Copyright 1991 by Analog Devices, Inc.
*
* Refer to "README.DOC" file for License Statement.  Use of this model
* indicates your acceptance with the terms and provisions in the License Statement.
*
* Node assignments
*              non-inverting input
*              | inverting input
*              | | positive supply
*              | | |   negative supply
*              | | |   |   output
*              | | |   |   |
.SUBCKT AD840J 1 2 100 101 36
*
* INPUT STAGE & POLE AT 120 MHz
*
IOS  1  2  DC  0.2E-6
CIN  1  2  2E-12
R1  1  3  3.2325E3
R2  2  3  3.2325E3
EOS  9  1  POLY(1)  16  11  1E-3  1
R3  100  5  195.45
R4  100  6  195.45
C2  5  6  3.3929E-12
R5  7  4  143.73
R6  8  4  143.73
Q1  5  2  7  QX
Q2  6  9  8  QX
I1  4  101  DC  1E-3
*
*  VIRTUAL NODE
*
RVN1  100  10  25E3
RVN2  10  101  25E3
*
* GAIN STAGE & DOMINANT POLE AT 3.8 KHz
*
EREF  11  0  10  0  1
G1  11  12  5  6  5.1163E-3
R7  12  11  14.659E6
C3  12  11  2.857E-12
V1  100  13  DC  5.0875
D1  12  13  DX
V2  14  101  DC  5.0875
D2  14  12  DX
*
* COMMON-MODE GAIN NETWORK WITH ZERO AT 200 KHz
*
ECM  15  11  3  11  31.623
RCM1  15  16  1E6
CCM  15  16  795.77E-15
RCM2  16  11  1
*
* NEGATIVE ZERO STAGE AT 290 MHz
*
EZ1  17  11  12  11  1E6
RZ1  17  18  1
CZ1  17  18  -548.81E-12
RZ2  18  11  1E-6
*
* POLE STAGE AT 500 MHz
*
GP1  11  19  18  11  1E-6
RP1  19  11  1E6
CP1  19  11  318.31E-18
*
* OUTPUT STAGE
*
IDC  100  101  DC  10.4E-3
VX  19  30
V3  32  35  DC  2.725
D3  30  32  DX
V4  35  33  DC  2.575
D4  33  30  DX
D5  100  31  DX
GO1  31  101  30  35  16.667E-3
D6  101  31  DY
D7  100  34  DX
GO2  34  101  35  30  16.667E-3
D8  101  34  DY
RO1  100  35  60
GO3  35  100  100  30  16.667E-3
RO2  35  101  60
GO4  101  35  30  101  16.667E-3
LO  35  36  0.04E-6
*
* MODELS USED
*
.MODEL QX NPN(BF=62.5)
.MODEL DX D(IS=1E-15)
.MODEL DY D(IS=1E-15 BV=50)
.ENDS
