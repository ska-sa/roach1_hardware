* ADG508F SPICE Macro-model                5/95, Rev. B
*                                          JOM / ADSC
*
* Revision History:
*     Rev A. S1-S8 label correction
*     Rev B. Leakage Currents
*     Rev C. Switching Times and Break before Make
*
*	NOTE: This model was setup with typical leakage currents
*		at +25 for ADG508F 
*
*        This model does not include the write and reset function.
*
* Copyright 1995 by Analog Devices, Inc.
*
* Refer to "README.DOC" file for License Statement.  Use of this 
* model indicates your acceptance with the terms and provisions 
* in the License Statement.
*
* Node assignments
* 4 - S1, 5 - S2, 6 - S3, 7 - S4, 12 - S5, 11 - S6, 10 - S7
* 9 - S8, 15 - A2, 16 - A1, 1 - A0, 2 - Enable, 8 - D
* 13 - Vdd, 14 - GND, 3 - Vss
*                    
.SUBCKT ADG508F 4 5 6 7 12 11 10 9 15 16 1 2 8 13 14 3
*
* DEMUX SWITCHES (S1-8 ---> D)
*
*     First Section is for control line A0
*          All nodes in this section are in the 30's unless
*          they are I/O nodes
*
E_A0_2	  200  0  1  0    1
E_A0_1     30 40 201 40   -1
R_A0_1    200 201         1000
C_A0_X2   201  0          130E-12

V_AX_1     40  0          1.6

S_A0_8      9 31 201 0	  Sdemux
S_A0_7     10 31 30  0	  Sdemux		
S_A0_6     11 32 201 0    Sdemux
S_A0_5     12 32 30  0    Sdemux
S_A0_4      7 33 201 0    Sdemux
S_A0_3      6 33 30  0    Sdemux
S_A0_2      5 34 201 0    Sdemux
S_A0_1      4 34 30  0    Sdemux

C_A0_X1     1  0          1E-12
C_A0_D      1 38          1E-12

*          Input capacitances

C_A0_1      4  0          5E-12
C_A0_2      5  0          5E-12
C_A0_3      6  0 	  5E-12
C_A0_4      7  0          5E-12
C_A0_5     12  0          5E-12
C_A0_6     11  0          5E-12
C_A0_7     10  0          5E-12
C_A0_8      9  0          5E-12

C_D_1       8  0          50E-12

*
*	Leakage Current (SX and D ON only) 
*

G_ON_S1     4  0  4  0    2E-12
G_ON_S2	    5  0  5  0    2E-12
G_ON_S3     6  0  6  0    2E-12
G_ON_S4     7  0  7  0    2E-12
G_ON_S5    12  0 12  0    2E-12
G_ON_S6    11  0 11  0    2E-12
G_ON_S7    10  0 10  0    2E-12
G_ON_S8     9  0  9  0    2E-12
G_ON_D	    8  0  8  0    2E-12		  

*
*	Leakage Current (SX OFF only
*
*	Leakage Current (D OFF only)
*

S_OFF_D     8  58 80  0	  Sdemux
R_OFF_D     58  0         1E12 
G_OFF_D     8   0 58  0   2E-12

*
*     Second Section is for control line A1
*

E_A1_2	  170  0 16  0    1
E_A1_1     37 40 171 40   -1
R_A1_1    170 171         1000
C_A1_X2   171  0          130E-12

S_A1_1     31 35 171 0     Sdemux
S_A1_2     32 35 37  0     Sdemux
S_A1_3     33 36 171 0     Sdemux
S_A1_4     34 36 37  0     Sdemux

C_A1_X     16  0           1E-12
C_A1_D     16 38           1E-12

*
*     Third Section is for control line A2
*

E_A2_2	  160  0 15  0    1
E_A2_1     39 40 161 40   -1
R_A2_1    160 161         1000
C_A2_X2   161  0          130E-12

S_A2_1     35 38 161 0     Sdemux
S_A2_2     36 38 39  0     Sdemux

C_A2_X     15  0           1E-12
C_A2_D     15 38           1E-12

*
*     Main Series Switch combination
*

S_1_E     41  73 611 0     SMAINP
S_1_F     380  41 612 0     SMAINN

E_1_E     611 0   VALUE = {(10*V(8,0))/(V(13,14)+0.15)}
E_1_F     612 0   VALUE = {(10*V(8,0))/(V(3,14)+0.15)}

SBASE     38  380  13  3  SBASE

*
*     Enable Switch section
*

S_EN_1     73  8  2  0     Sdemux
C_EN_1      2 73           3E-12

*     Invert Enable Switch section

E_EN0_1     80  0  2  81   -2
V_EN0_1	    81  0          2.5

*
*     Power Supply Current Correction
*
I_PS_1     13  0           0.05E-3
I_PS_2      0  3           0.01E-3
E_PS_1     99  0 13  0     1

*
* MODELS USED
*
.MODEL SBASE  VSWITCH(RON=260 ROFF=1200 VON=30 VOFF=-10)
.MODEL SMAINN VSWITCH(RON=10000 ROFF=3 VON=13 VOFF=0)
.MODEL SMAINP VSWITCH(RON=10000 ROFF=3 VON=13 VOFF=0)
.MODEL Sdemux VSWITCH (RON=1 ROFF=1E12 VON=2.0 VOFF=1.4)
.ENDS ADG508F
