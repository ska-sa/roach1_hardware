* ADG426 SPICE Macro-model                10/95, Rev. D
*                                           WF / ADSC
*
* Revision History: NONE
*
*       NOTES: 1. This model was setup with typical leakage currents
*               at +25C for ADG426 
*              2. The digital address latches are not implemented.
*
* Copyright 1995 by Analog Devices, Inc.
*
* Refer to "README.DOC" file for License Statement.  Use of this 
* model indicates your acceptance with the terms and provisions 
* in the License Statement.
*
* Node assignments
* 19 - S1, 20 - S2, 21 - S3, 22 - S4, 23 - S5, 24 - S6, 25 - S7
* 26 - S8, 11 - S9,10 - S10, 9 - S11, 8 - S12, 7 - S13, 6 - S14
* 5 - S15, 4 - S16, 14 - A3, 15 - A2, 16 - A1, 17 - A0, 18 - EN
* 28 - D, 1 - VDD, 12 - GND, 27 - VSS
*                    
.SUBCKT ADG426 19 20 21 22 23 24 25 26 11 10 9 8 7 6 5 4 14 15 16 17 18 28 1 12 27
*
* DEMUX SWITCHES (S1-16 ---> D)
*
*     First Section is for control line A0
*          All nodes in this section are in the 30's unless
*          they are I/O nodes
*
E_A0_2    200 12  17 12    1
E_A0_1     30 40 201 40   -1
R_A0_1    200 201         1000
C_A0_X2   201 12          100E-12

V_AX_1     40  12          1.6

S_A0_16     4 31 201 12   Sdemux
S_A0_15     5 31 30  12   Sdemux                
S_A0_14     6 32 201 12   Sdemux
S_A0_13     7 32 30  12   Sdemux
S_A0_12     8 33 201 12   Sdemux
S_A0_11     9 33 30  12   Sdemux
S_A0_10    10 34 201 12   Sdemux
S_A0_9     11 34 30  12   Sdemux
S_A0_8     26 35 201 12   Sdemux
S_A0_7     25 35 30  12   Sdemux                
S_A0_6     24 36 201 12   Sdemux
S_A0_5     23 36 30  12   Sdemux
S_A0_4     22 37 201 12   Sdemux
S_A0_3     21 37 30  12   Sdemux
S_A0_2     20 38 201 12   Sdemux
S_A0_1     19 38 30  12   Sdemux

C_A0_X1     17 12          4E-12
C_A0_D      17 39          4E-12

*          Input capacitances

C_A0_1     19  12          8E-12
C_A0_2     20  12         8E-12
C_A0_3     21  12         8E-12
C_A0_4     22  12         8E-12
C_A0_5     23  12         8E-12
C_A0_6     24  12         8E-12
C_A0_7     25  12         8E-12
C_A0_8     26  12         8E-12
C_A0_9     11  12         8E-12
C_A0_10    10  12         8E-12
C_A0_11     9  12         8E-12
C_A0_12     8  12         8E-12
C_A0_13     7  12         8E-12
C_A0_14     6  12         8E-12
C_A0_15     5  12         8E-12
C_A0_16     4  12         8E-12

C_D_1      28  12         80E-12

*
*       Leakage Current (SX and D ON only) 
*

R_ON_S1    19 500    1.5E12
R_ON_S2    20 500    1.5E12
R_ON_S3    21 500    1.5E12
R_ON_S4    22 500    1.5E12
R_ON_S5    23 500    1.5E12
R_ON_S6    24 500    1.5E12
R_ON_S7    25 500    1.5E12
R_ON_S8    26 500    1.5E12
R_ON_S9    11 500    1.5E12
R_ON_S10   10 500    1.5E12
R_ON_S11    9 500    1.5E12
R_ON_S12    8 500    1.5E12
R_ON_S13    7 500    1.5E12
R_ON_S14    6 500    1.5E12
R_ON_S15    5 500    1.5E12
R_ON_S16    4 500    1.5E12
SLEAK_ON_D 28 500    28 500  SLEAK
ILEAK_ON_D 28 500   -10E-12               
* 
*       Leakage Current (SX OFF only)
*
*       Leakage Current (D OFF only)
*
S_OFF_D     28  58 80 12          Sdemux
R_OFF_D     58  12                1E12 
G_OFF_D     28  12 58 12          0.75E-12
*
*     Second Section is for control line A1
*
E_A1_2    170 12 16  12    1
E_A1_1     41 40 171 40   -1
R_A1_1    170 171         1000
C_A1_X2   171 12          100E-12
*
S_A1_1     31 42 171 12     Sdemux
S_A1_2     32 42 41  12     Sdemux
S_A1_3     33 43 171 12    Sdemux
S_A1_4     34 43 41  12    Sdemux
S_A1_5     35 44 171 12    Sdemux
S_A1_6     36 44 41  12    Sdemux
S_A1_7     37 45 171 12    Sdemux
S_A1_8     38 45 41  12    Sdemux
*
C_A1_X     16 12           4E-12
C_A1_D     16 39           4E-12
*
*     Third Section is for control line A2
*

E_A2_2    160 12 15  12    1
E_A2_1     46 40 161 40   -1
R_A2_1    160 161         1000
C_A2_X2   161  12          100E-12

S_A2_1     42 47 161 12     Sdemux
S_A2_2     43 47 46  12    Sdemux
S_A2_3     44 48 161 12    Sdemux
S_A2_4     45 48 46  12    Sdemux

C_A2_X     15 12           4E-12
C_A2_D     15 39           4E-12

*
*     Forth Section is for control line A3
*

E_A3_2    140  12  14 12   1
E_A3_1     49  40 141 40   -1
R_A3_1    140 141         1000
C_A3_X2   141  12          100E-12

S_A3_1     47 39 141 12     Sdemux
S_A3_2     48 39 49  12    Sdemux

C_A3_X     14 12           4E-12
C_A3_D     14 39           4E-12

*
*     Main Series Switch combination
*
*

V_1_A     419  12  15
V_1_B     420  12  -15
V_1_C     421  500 -0.5         ;sets pos main offset
V_1_D     422  27  2.5          ;sets neg main offset
R_1_C     39   0   1E13
S_1_A     425  39  420 73 SNCM
R_1_A    412 425  24            ;sets neg at max d
S_1_B      426  39  419 73 SPCM
R_1_B     73 426  30            ;sets pos at max d
S_1_C      73 412 611  12 SMAINP
S_1_D     412 411  12 612 SMAINN
E_1_E     611  12         VALUE = {(10*V(73,421))/(0.5*V(1,500)+0.005)}
E_1_F     612  12         VALUE = {(10*V(73,500))/(PWR(V(500,422),1)+0.005)}
S_1_G     411  39   1  27 SBASE

I_XX_1    99 0 0       ;add a 'do-nothing' component
I_XX_3   421 0 0      ;  at nodes 99, 421
I_XX_3   422 0 0      ;    and 422 to keep SPICE happy

*
*       Voltage Clamp 
*

D_1_POS     39  1    DClamp
G_1_POS     39  1  39  1  -1E-12
D_2_NEG     27  39   DClamp
G_2_NEG     27  39 27  39 1E-12

*     Enable Switch section
*

S_EN_1     73 28 18  12     Sdemux
C_EN_1     18 28           4.2E-12  ; SETS CHARGE INJECTION 

*     Invert Enable Switch section

E_EN0_1     18  81 80 12    -2
V_EN0_1     82  12          2.5
R_EN0_1     82  81         1
R_EN0_2     80  12          1E12

*
*     Power Supply Current Correction
*
I_PS_1      1  12           80E-6
I_PS_2     12  27           0.0001E-6
E_PS_1     99  12  1  12    1
E_PS_2    500  27  1  27    .5

*
*       Crosstalk 
*

RXT_1     19 52           1E13
RXT_2     20 52           1E13
RXT_3     21 52           1E13
RXT_4     22 52           1E13
RXT_5     23 52           1E13
RXT_6     24 52           1E13
RXT_7     25 52           1E13
RXT_8     26 52           1E13
RXT_9     11 52           1E13
RXT_10    10 52           1E13
RXT_11     9 52           1E13
RXT_12     8 52           1E13
RXT_13     7 52           1E13
RXT_14     6 52           1E13
RXT_15     5 52           1E13
RXT_16     4 52           1E13

CXT_1     19 52           1E-12
CXT_2     20 52           1E-12
CXT_3     21 52           1E-12
CXT_4     22 52           1E-12
CXT_5     23 52           1E-12
CXT_6     24 52           1E-12
CXT_7     25 52           1E-12
CXT_8     26 52           1E-12
CXT_9     11 52           1E-12
CXT_10    10 52           1E-12
CXT_11     9 52           1E-12
CXT_12     8 52           1E-12
CXT_13     7 52           1E-12
CXT_14     6 52           1E-12
CXT_15     5 52           1E-12
CXT_16     4 52           1E-12

*
*       OFF Isolation
*
COI_1     19 28           1E-13
COI_2     20 28           1E-13
COI_3     21 28           1E-13
COI_4     22 28           1E-13
COI_5     23 28           1E-13
COI_6     24 28           1E-13
COI_7     25 28           1E-13
COI_8     26 28           1E-13
COI_9     11 28           1E-13
COI_10    10 28           1E-13
COI_11     9 28           1E-13
COI_12     8 28           1E-13
COI_13     7 28           1E-13
COI_14     6 28           1E-13
COI_15     5 28           1E-13
COI_16     4 28           1E-13
ROI_1     19 1901         1.6E9
COI_1A    1901 28         10E-12
ROI_2     20 1902         1.6E9
COI_2A    1902 28         10E-12
ROI_3     21 1903         1.6E9
COI_3A    1903 28         10E-12
ROI_4     22 1904         1.6E9
COI_4A    1904 28         10E-12
ROI_5     23 1905         1.6E9
COI_5A    1905 28         10E-12
ROI_6     24 1906         1.6E9
COI_6A    1906 28         10E-12
ROI_7     25 1907         1.6E9
COI_7A    1907 28         10E-12
ROI_8     26 1908         1.6E9
COI_8A    1908 28         10E-12
ROI_9     11 1909         1.6E9
COI_9A    1909 28         10E-12
ROI_10     10 1910         1.6E9
COI_10A    1910 28         10E-12
ROI_11     9 1911         1.6E9
COI_11A    1911 28         10E-12
ROI_12     8 1912         1.6E9
COI_12A    1912 28         10E-12
ROI_13     7 1913         1.6E9
COI_13A    1913 28         10E-12
ROI_14     6 1914         1.6E9
COI_14A    1914 28         10E-12
ROI_15     5 1915         1.6E9
COI_15A    1915 28         10E-12
ROI_16     4 1916         1.6E9
COI_16A    1916 28         10E-12
*
* MODELS USED
*
.MODEL SNCM  VSWITCH (RON=1 ROFF=500001 VON=9 VOFF=-44)
.MODEL SPCM  VSWITCH (RON=450000 ROFF=1 VON=41 VOFF=-6.5)
.MODEL SBASE VSWITCH (RON=11 ROFF=3500 VON=28 VOFF=-10)
.MODEL SMAINP VSWITCH (RON=650001 ROFF=19 VON=32 VOFF=0)
.MODEL SMAINN VSWITCH (RON=700001 ROFF=7 VON=28.5 VOFF=0)
.MODEL Sdemux VSWITCH (RON=1 ROFF=1E12 VON=2.0 VOFF=1.4)
.MODEL DClamp D(IS=1E-15 IBV=1E-13)
.MODEL SLEAK VSWITCH (RON=750E9 ROFF=150E9 VON=-15 VOFF=15)
.ENDS ADG426
