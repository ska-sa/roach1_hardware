* ADN8830 Mixed Signal SPICE Model v0.2
*
* Copyright 2001 Analog Devices, Inc.
* TAM 11/01
*
* Note: Node numbers 1-32 refer to actual pin numbers on device
*
.SUBCKT ADN8830_M 1 2 3 4 5 6 7 8 9 10 11 12 13 14 17 18 19
+ 20 21 22 23 24 25 26 27 28 29 30 31 
*
* CLOCK SECTION
*
V15    6 30 1.5V
V30   33 30 3V
VFREQ 26 30 3V
F1 30 66 POLY(2) V5 VFREQ 0 0 0 0 100E3
C1 66 30 333p     ; with I(VFREQ)=20uA, dV/dt=6V/1us
R3 66 30 100E3  ; 100E6

O1 66 33 ADCONV DGTLNET=50 IO_CMOS
O2 30 66 ADCONV DGTLNET=51 IO_CMOS
U7 SRFF(1) 8 30 DIG1 DIG1 DIG1
+          50 51 52 53 T_SRF IO_CMOS ; 52 is Q output
U10 PULLUP(1) 8 30 DIG1 R1K

N3 60 30 33 DACONV DGTLNET=52 IO_CMOS
R1 60 61 1.5k
V5 61 30 1.5V ; current through V1 should be +1mA or -1mA
N4 28 30  8 DACONV DGTLNET=52 IO_CMOS
*
* PWM Duty Cycle Control
*
O3 17 66 ADCONV  DGTLNET=42       IO_CMOS
U1 INV     20 23 42 43    T_STD   IO_CMOS
U2 DLYLINE 20 23 43 44    DLY80NS IO_CMOS
U3 NAND(2) 20 23 43 44 45 T_STD   IO_CMOS
U4 INV     20 23 44 46    T_STD   IO_CMOS
U5 NAND(2) 20 23 42 46 47 T_STD   IO_CMOS
U6 INV     20 23 45 48    T_STD   IO_CMOS
N1 22 23 20 DACONV DGTLNET=48     IO_CMOS
N2 21 23 20 DACONV DGTLNET=47     IO_CMOS
*
* THERMFAULT Output
*
V6 71 30 2.3V
V7 72 30 0.2V
O4  2 71 ADCONV  DGTLNET=54  IO_CMOS
O5 72  2 ADCONV  DGTLNET=55  IO_CMOS
U8 OR(2) 8 30 54 55 56 T_STD IO_CMOS
N5  1 30 8 DACONV DGTLNET=56 IO_CMOS
*
* TEMPLOCK Output
*
V8 73 30 1.55V
V9 74 30 1.45V
O6 73 12 ADCONV DGTLNET=57    IO_CMOS
O7 12 74 ADCONV DGTLNET=58    IO_CMOS
U9 AND(2) 8 30 57 58 59 T_STD IO_CMOS
N6  5 30  8 DACONV DGTLNET=59 IO_CMOS
*
* Linear Output Amplifier
*
R2  14 89 10k
R4  89  9 140k
G1  20 11 (89,6) 37.7m
R19 11 20 147.4k
D1  11 85 DX
V1  20 85 0.75
D2  86 11 DX
V2  86 23 0.75
G2  23 10 (89,6) 37.7m
R20 10 23 603.2k
D3  10 87 DX
V3  20 87 0.75
D4  88 10 DX
V4  88 23 0.75
*
* PWM Control Voltage Section
*
E1  80 30 POLY(2) (14,30) (9,30) 9 -4 -1
R17 80 18 100k
R18 18 19 100k
X1   6 18 17 33 30 OPAMP
*
* Compensation Amplifier
*
X2   6 13 14 33 30 OPAMP
*
* Input Error Amplifier
*
E2  34  6 POLY(1) (4,2) 0 20 ; (TEMPSET-THERMIN)*20 + 1.5V
R9  34 12 0.1
VREF 7 30 2.45V
*
* TEMPOUT Amplifier
*
E3  35  6 (4,2) 3
R10 35 31 0.1
*
* Dummy Pins
*
RSY  8 30 100k ; AVDD to AGND ISY
* R32 32 30 1MEG
R25 25 30 1MEG
R29 29 30 1MEG
R24  8 24 1k
R27 27 30 1MEG
RSD  3 30 1MEG
*
.MODEL ADCONV DOUTPUT(RLOAD=1E8,S0NAME="0",S0VLO=-5E4,S0VHI=0,
+                               S1NAME="1",S1VLO=0,S1VHI=5E4)
.MODEL T_STD UGATE()
.MODEL T_SRF UGFF()
.MODEL DLY80NS UDLY(DLYTY=80ns)
.MODEL DACONV DINPUT(S0NAME="0",S0TSW=20ns,S0RLO=2,S0RHI=5E6,
+                    S1NAME="1",S1TSW=20ns,S1RLO=5E6,S1RHI=2,
+                    S2NAME="X",S2TSW=20ns,S2RLO=5E6,S2RHI=5E6,
+                    S3NAME="Z",S3TSW= 1ns,S3RLO=5E6,S3RHI=5E6)
.MODEL IO_CMOS UIO()
.MODEL R1K UIO(DRVZ=1k,INR=30k)
* .MODEL NLINFET NMOS(LEVEL=2,KP=24E-6,VTO=1, LAMBDA=0.01)
* .MODEL PLINFET PMOS(LEVEL=2,KP=24E-6,VTO=-1,LAMBDA=0.01)
.MODEL DX D(IS=1E-14,RS=1m)
.ENDS
*
* Simple Op Amp Avo=120k
*
.SUBCKT OPAMP 1 2 3 99 50
G1 50  4 (2,1) 1
R1  4 50 100k
C1  4 50 1.5p
D1  4 98 DX
V1 99 98 0.6
D2 51  4 DX
V2 51 50 0.6
M1  3  4 50 50 NAMPFET L=1u W=10m
R2 99  3 10k
.MODEL DX D(IS=1E-14,RS=1m)
.MODEL NAMPFET NMOS(LEVEL=1,VTO=0,KP=24E-6)
.ENDS
*$