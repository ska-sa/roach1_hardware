* AD813A SPICE Macro-model                  11/93, Rev. A   
*                                           JCB / PMI
*
* This version of the AD813 model simulates the worst case 
* parameters of the 'A' grade.  The worst case parameters
* used correspond to those in the data sheet.  This model was
* developed using the +-5V specifications.
*
* Copyright 1993 by Analog Devices, Inc.
*
* Refer to "README.DOC" file for License Statement.
* Use of this model indicates your acceptance with
* the terms and provisions in the License Statement.
*
* Node assignments
*              non-inverting input
*              | inverting input
*              | | positive supply
*              | | |  negative supply
*              | | |  |  output
*              | | |  |  |  DISABLE pin
*              | | |  |  |  |     
.SUBCKT AD813A 1 2 99 50 41 33
*
* INPUT STAGE
*
R1   99  8     1000
R2   10 50     1000
V1   99  9     -0.15
D1   9   8     DX
V2   11 50     -0.15
D2   10 11     DX
F1   99  5     VD2  1
F2   4  50     VD2  1
Q1   50  3  5  QP
Q2   99  3  4  QN
Q3   8   5  2  QN
Q4   10  4  2  QP
R3   99  5     0.4E8
R4   50  4     0.4E8
*
* INPUT ERROR SOURCES
* 
GB1  99  1     POLY(1)  1  22  1.5E-6  150E-9
GB2  99  2     POLY(1)  1  22  30E-6  3E-6
EOS  3   1     POLY(1)  16 22  5E-3  1
CS1  99  2     0.75E-12
CS2  99  1     1.7E-12
*
EREF 97  0     22  0  1
*
* TRANSCONDUCTANCE STAGE
*
R5   12 97     1.2E6
C3   12 97     4.3E-12
G1   97 12     99  8  1E-3
G2   12 97     10 50  1E-3
V3   99 13     1.85
V4   14 50     1.85
D3   12 13     DX
D4   14 12     DX
*
* COMMON-MODE GAIN NETWORK WITH ZERO AT 19 KHZ
*
R11  15 16   1E4
R12  16 97   1
C5   15 16   5E-12
E3   97 15   1  22  12
*
* POLE AT 100 MHZ
*
R6   21 97    1E6
C4   21 97    1.59E-15
G3   97 21    12 22  1E-6
*
* OUTPUT STAGE
*
FSY  99 50    POLY(1)  VD2  0.5E-3  14
FSY1 99  0    V7  1
FSY2 0  50    V8  1
R9   22 99    10E3
R10  22 50    10E3
E1   25 97    21 22 1
H1   26 25    POLY(1) VD3 0.68 10E3
H2   25 27    POLY(1) VD3 0.68 10E3
RH1  40 50    1E10
R7   28 40    10
R8   40 29    10
D7   26 28    DX
D8   29 27    DX
VS   40 41    DC 0
CL   41 50    10E-12
V5   23 40    0.55
V6   40 24    0.55
D5   21 23    DX
D6   24 21    DX
*
F10  97 70    VS 1
D9   70 71    DX
D10  72 70    DX
V7   71 97    DC 0
V8   97 72    DC 0
*
* DISABLE FUNCTION
*
VD1  99 31    DC 1.8
RD1  31 32    35E3
RD2  33 99    1E12
DD1  32 33    DX
FD   97 34    POLY(1) VD1 215E-6 -10
DD3  36 34    DX
DD2  34 35    DX
VD2  37 97    DC 0
VD3  38 97    DC 0
RD3  35 37    1E3
RD4  36 38    1E3
CD1  34 97    10E-12
*
* MODELS USED
*
.MODEL QN   NPN(BF=200 IS=1E-15)
.MODEL QP   PNP(BF=200 IS=1E-15)
.MODEL DX   D(IS=1E-15)
.ENDS
