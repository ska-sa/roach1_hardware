* AD8210 SPICE Macro-Model	REV 0, 3/2006, TRW, ADI
*
* Refer to "README.DOC" file for License Statement.
* Use of this model indicates your acceptance with
* the terms and provisions in the License Statement.
*
* The following parameters are accurately modeled;
*
*       Closed loop gain vs. frequency
*       output impedance 
*       output clamping voltage and current
*       CMRR
*       slew rate
*       distortion is not characterized       
*
*
*    Node assignments
*              non-inverting input
*              | inverting input
*              | |  positive supply
*              | |  |  negative supply
*              | |  |  |  Vref+
*              | |  |  |  |  Vref-
*              | |  |  |  |  | output
*              | |  |  |  |  | |

.subckt AD8210 1 83 99 50 8 9 45

*** Reference Stage

Eref 98 0 poly(2) 99 0 50 0 0 0.5 0.5
Erefout 97 0 poly(2) 8 0 9 0 0 0.5 0.5
Iq 50 99 24.996

*** Input Stage

Eos 83 2 poly(1) 66 98 0 .05 
*Vos 83 2 0
Vref+ 9999 0 65
Vref- 0 5000 2
Eref+ 999 0 9999 0 1
Eref- 0 500 0 5000 2
Ecm 65 0 poly(2) 1 0 2 0 0 0.5 0.5
Rcm1 65 66 1meg
Rcm2 66 98 1
Ccm 65 66 79p

Rindiff 1 2 2k
Rincm1 1 98 10Meg
Rincm2 2 98 10Meg

Q1 4 1 5 NPN
Q2 3 2 6 NPN
I1 7 500 1
Rc1 999 3 50
Rc2 999 4 50
Re1 5 7 49
Re2 6 7 49

*** Gain Stage

Gd1 13 98 4 3 20.894
Rd1 13 98 0.955
Cd1 13 98 3.33e-7

*** Output clamping

D1 13 14 dx
D2 15 13 dx
Vd1 14 99 -1.025
Vd2 15 50 0.87

Ebuf 97 21 13 98 1
Gbuf 22 98 21 97 .01
Rbuf 98 22 100
Dout1 23 22 dx
Dout2 22 24 dx
Vout1 45 23 -.6
Vout2 24 45 -.6

Gout1 45 99 98 22 .5
Gout2 50 45 22 98 .5
Rout1 45 99 2
Rout2 50 45 2

.model npn npn(bf=2500)
.model dx D
.ends
