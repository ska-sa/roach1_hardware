* AD843J  SPICE Macro-model                 1/92, Rev. A
*                                           JCB / PMI
*
* This version of the AD843 model simulates the worst case 
* parameters of the 'J' grade.  The worst case parameters
* used correspond to those in the data sheet.
*
* Copyright 1991 by Analog Devices, Inc.
*
* Refer to "README.DOC" file for License Statement.  Use of this model
* indicates your acceptance with the terms and provisions in the License Statement.
*
* Node assignments
*                non-inverting input
*                | inverting input
*                | | positive supply
*                | | |  negative supply
*                | | |  |  output
*                | | |  |  |
.SUBCKT AD843J   1 2 99 50 30
*
* INPUT STAGE & POLE AT 150 MHZ
*
R1   1   3   5E11
R2   2   3   5E11
R3   5  50   693.9
R4   6  50   693.9
CIN  1   2   4E-12
C2   5   6   0.765E-12
I1   99  4   1.0E-3
IOS  1   2   5E-10
EOS  7   1   POLY(1)  16 24  2E-3  1
J1   5   2   4   JX
J2   6   7   4   JX
*
EREF 98  0   24  0  1
*
* GAIN STAGE & POLE AT 2.45 KHZ
*
R5   9  98   1.04E7
C3   9  98   6.25E-12
G1   98  9   5  6  1.44E-3
V2   99  8   5.2
V3   10 50   5.2
D1   9   8   DX
D2   10  9   DX
*
* POLE AT 200 MHZ
*
R6   11 98   1E6
C4   11 98   0.796E-15
G2   98 11   9 24  1E-6
*
* NEGATIVE ZERO AT 100 MHZ
*
R8   13 14   1E6
R9   14 98   1
C6   13 14   -1.59E-15
E2   13 98   11  24  1000001
*
* COMMON-MODE GAIN NETWORK WITH ZERO AT 120 KHZ
*
R10  15 16   1E6
R11  16 98   1
C7   15 16   1.326E-12
E3   98 15   3  24  1000
*
* POLE AT 200 MHZ
*
R12  23 98   1E6
C8   23 98   0.796E-15
G4   98 23   14  24  1E-6
*
* OUTPUT STAGE
*
R13  24 99   50E3
R14  24 50   50E3
ISY  99 50   11.7E-3
R15  29 99   40
R16  29 50   40
L1   29 30   6E-8
G5   27 50   23 29  2.5E-2
G6   28 50   29 23  2.5E-2
G7   29 99   99 23  2.5E-2
G8   50 29   23 50  2.5E-2
V4   25 29   0.3
V5   29 26   0.3
D3   23 25   DX
D4   26 23   DX
D5   99 27   DX
D6   99 28   DX
D7   50 27   DY
D8   50 28   DY
*
* MODELS USED
*
.MODEL JX PJF(BETA=1.04E-3  VTO=-2.000  IS=2.5E-9)
.MODEL DX   D(IS=1E-15)
.MODEL DY   D(IS=1E-15 BV=50)
.ENDS
