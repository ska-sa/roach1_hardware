* OP193E SPICE Macro-model              1/95, Rev. A
*                                       ARG / ADI
*
* This version of the OP193 model simulates the worst-case
* parameters of the 'E' grade.  The worst-case parameters
* used correspond to those in the data sheet.
*
* Copyright 1990 by Analog Devices, Inc.
*
* Refer to "README.DOC" file for License Statement. Use of this model
* indicates your acceptance with the terms and provisions in the License
* Statement. This model has been optimized for a total supply voltage of
* 5V.
*
* Node assignments
*              non-inverting input
*              |  inverting input
*              |  |  positive supply
*              |  |  |  negative supply
*              |  |  |  |  output
*              |  |  |  |  |
.SUBCKT OP193E 51 52 99 50 32
*
* INPUT STAGE & POLE AT 16KHZ
*
R3   5    50   53.827E3
R4   6    50   53.827E3
R5   4    7    2.104E3
R6   4    8    2.104E3
CIN  1    2    4E-12
C2   5    6    92.4E-12
I1   99   4    1.03E-6
IOS  1    2    1E-9
EOS  9    1    POLY(2) (24,27) (102,0) 75E-6 0.1 1
Q1   5    2    7    QX
Q2   6    9    8    QX
EREF 98   0    POLY(2) (99,0) (50,0) 0 0.5 0.5
R24  1    51   2E3
R25  2    52   2E3
VN1  101  0    DC 2
VN2  0    103  DC 2
DN1  101  102  DEN
DN2  102  103  DEN
*
* GAIN STAGE & DOMINANT POLE AT 0.473 HZ
*
R7   10   98   4.037E9
G1   98   10   (5,6) 18.578E-6
C3   10   98   83.333E-12
V1   99   11   0.65
D1   10   11   DX
D2   50   10   DX
*
* NEGATIVE ZERO AT 50KHZ
*
R9   13   14   1E6
R10  14   98   1
FNZ  13   14   VNZ -1
E2   13   98   (10,27) 1
CNZ  15   16   3.183E-12
ENZ  15   98   (13,14) 1
VNZ  16   98   DC 0
*
* ZERO-POLE PAIR AT 28KHZ / 84KHZ
*
R18  17   18   2E6
C4   17   18   2.842E-12
R19  18   98   1E6
E3   17   98   (14,27) 3E6
*
* COMMON-MODE GAIN NETWORK WITH ZERO AT 3.16HZ
*
R1   23   24   1E6
R2   24   98   100
C5   23   24   50.33E-9
E4   23   98   POLY(2) (1,27) (2,27) 0 0.5 0.5
*
* ZERO-POLE PAIR AT 40KHZ / 160KHZ
*
R20  25   26   3E6
C6   25   26   1.326E-12
R21  26   98   1E6
E5   25   98   (18,27) 4
*
* OUTPUT STAGE
*
ISY  99   50   20.137E-6
R16  27   99   4.5E6
R17  27   50   4.5E6
EIN  28   98   POLY(1) (26,27) 0.51905 1
RIN  28   31   15E3
Q11  45   31   32   QN 6
Q12  32   33   44   QN 6
Q13  41   34   33   QN 1
Q14  34   35   36   QP 1
Q15  36   38   39   QN 8
Q16  35   35   37   QP 1
Q17  99   99   37   QN 1
Q18  99   99   36   QN 1
Q19  50   42   34   QP 1
Q20  42   42   34   QP 1
Q21  32   33   42   QN 1
Q22  99   40   41   QN 1
Q23  43   43   50   QN 1
Q24  34   43   50   QN 2
Q25  33   43   50   QN 2
Q26  34   44   50   QC 1
Q27  31   46   50   QC 1
EC   47   50   (99,45) 0.96
RC   46   47   1E3
IREF 99   43   4.5E-7
I13  35   50   4.5E-7
R11  99   40   75E3
R12  99   36   40E3
R13  31   38   20E3
R14  32   39   5E3
R15  40   37   75E3
R22  44   50   30
R23  99   45   50
*
* MODELS USED
*
.MODEL QN NPN(BF=200 IS=1E-16 VA=150)
.MODEL QP PNP(BF=100 IS=5E-17 VA=50)
.MODEL QX PNP(BF=33.333 KF=2E-17)
.MODEL QC NPN(BF=200 IS=2.22E-11)
.MODEL DX D(IS=1E-15)
.MODEL DEN D(RS=2.45E3 KF=33E-15)
.ENDS
