* AD812 SPICE Macro-model                   12/93, Rev. A   
*                                           JCB / PMI
*
* Copyright 1993 by Analog Devices, Inc.
*
* This model was developed using the +-5V specifications.
*
* Refer to "README.DOC" file for License Statement.
* Use of this model indicates your acceptance with
* the terms and provisions in the License Statement.
*
* Node assignments
*              non-inverting input
*              | inverting input
*              | | positive supply
*              | | |  negative supply
*              | | |  |  output
*              | | |  |  |
.SUBCKT AD812  1 2 99 50 28
*
* INPUT STAGE
*
R1   99  8     1E3
R2   10 50     1E3
V1   99  9     1.3
D1   9   8     DX
V2   11 50     1.3
D2   10 11     DX
I1   99  5     140E-6
I2   4  50     140E-6
Q1   5   5  3  QN
Q2   4   4  3  QP
Q3   8   5  2  QN
Q4   10  4  2  QP
*
* INPUT ERROR SOURCES
* 
GB1  99  1     POLY(1)  1  22  0.3E-6  0.07E-6
GB2  99  2     POLY(1)  1  22  7E-6  2E-6
EOS  3   1     POLY(1)  16 22  2E-3  1
CS2  50  2     1.7E-12
CIN  1  50     1.7E-12
*
EREF 98  0     22  0  1
*
* GAIN STAGE & DOMINANT POLE
*
R5   12 98     1.2E6
C3   12 98     3.8E-12
G1   98 12     99  8  1E-3
G2   12 98     10 50  1E-3
V3   99 13     1.1
V4   14 50     1.1
D3   12 13     DX
D4   14 12     DX
*
* POLE AT 200 MHZ
*
R6  17 98     1E6
C4  17 98     0.795E-15
G3  98 17     12 22  1E-6
*
* COMMON-MODE GAIN NETWORK WITH ZERO AT 19 KHZ
*
R7  15 16   1E4
R8  16 98   1
C5  15 16   30E-12
E3  98 15   1  22  7.0
*
* POLE AT 150 MHZ
*
R9  21 98     1E6
C6  21 98     1.06E-15
G4  98 21     17 22  1E-6
*
* OUTPUT STAGE
*
R10 22 99     8E3
R11 22 50     8E3
R12 27 99     60
R13 27 50     60
L2  27 28     1E-8
G5  27 99     99 21  16.67E-3
G6  50 27     21 50  16.67E-3
V5  23 27     1.75
V6  27 24     1.75
D5  21 23     DX
D6  24 21     DX
G7  98 35     (27,21)  16.67E-3
D7  35 36     DX
D8  37 35     DX
V7  36 98     DC 0
V8  98 37     DC 0
F1  99 50     POLY(2) V7 V8 2.604E-3  1  1
*
* MODELS USED
*
.MODEL QN   NPN(BF=1E3 IS=1E-15)
.MODEL QP   PNP(BF=1E3 IS=1E-15)
.MODEL DX   D(IS=1E-15)
.ENDS
