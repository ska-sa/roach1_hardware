* Netlist for net Lsw00 - C:\Work\Roach\elec\SISim\PPC_DDR2\_1I289_PPC_ECC6.sp


* Output from HyperLynx SPICE Writer
* Created by . on Date: Monday Mar. 3,2008   Time: 8:26:58
* Created with HyperLynx version: 7.7 build: 385
* Design file: $1I289_PPC_ECC6.ffs
* Special Settings: Coupled


.SUBCKT _1I289_PPC_ECC6 Vinp Vinn 101 106 108 104 105 114 120 303 126 304 132 305 138 306 144 307 150 308 156 309
+  162 310 168 311 174 312 180 313 186 314 192 315 198 316 204 317 210 318 216 319
+  222 320 228 321 234 322 240 323 246 324 252 325 258 326 264 327 270 328 276 329
+  282 330 288 331 294 332 296 301

* Node  #  = <Reference Designator>.<pin name>
**********************************************
* Node 101 = EBD-J8_C249.1 (at pin)
* Node 106 = EBD-J8_R102.2 (at pin)
* Node 108 = EBD-J8_R102.1 (at pin)
* Node 104 = EBD-J8_U15.J9 (at pin) (receiver)
X_mdl_109 109 d_receive_109 MODEL_EBD-J8_U15_J9_ip
* Node 105 = EBD-J8_U5.J1 (at pin) (receiver)
X_mdl_111 111 d_receive_111 MODEL_EBD-J8_U5_J1_ip
* Node 114 = J10.17 (at pin)
* Node 120 = J10.32 (at pin)
* Node 303 = R32.2 (at pin)
* Node 126 = J10.31 (at pin)
* Node 304 = R31.2 (at pin)
* Node 132 = J10.30 (at pin)
* Node 305 = R30.2 (at pin)
* Node 138 = J10.29 (at pin)
* Node 306 = R29.2 (at pin)
* Node 144 = J10.28 (at pin)
* Node 307 = R28.2 (at pin)
* Node 150 = J10.27 (at pin)
* Node 308 = R27.2 (at pin)
* Node 156 = J10.26 (at pin)
* Node 309 = R26.2 (at pin)
* Node 162 = J10.25 (at pin)
* Node 310 = R25.2 (at pin)
* Node 168 = J10.24 (at pin)
* Node 311 = R24.2 (at pin)
* Node 174 = J10.23 (at pin)
* Node 312 = R23.2 (at pin)
* Node 180 = J10.22 (at pin)
* Node 313 = R22.2 (at pin)
* Node 186 = J10.21 (at pin)
* Node 314 = R21.2 (at pin)
* Node 192 = J10.20 (at pin)
* Node 315 = R20.2 (at pin)
* Node 198 = J10.19 (at pin)
* Node 316 = R19.2 (at pin)
* Node 204 = J10.18 (at pin)
* Node 317 = R18.2 (at pin)
* Node 210 = J10.16 (at pin)
* Node 318 = R16.2 (at pin)
* Node 216 = J10.15 (at pin)
* Node 319 = R15.2 (at pin)
* Node 222 = J10.14 (at pin)
* Node 320 = R14.2 (at pin)
* Node 228 = J10.13 (at pin)
* Node 321 = R13.2 (at pin)
* Node 234 = J10.12 (at pin)
* Node 322 = R12.2 (at pin)
* Node 240 = J10.11 (at pin)
* Node 323 = R11.2 (at pin)
* Node 246 = J10.10 (at pin)
* Node 324 = R10.2 (at pin)
* Node 252 = J10.9 (at pin)
* Node 325 = R9.2 (at pin)
* Node 258 = J10.8 (at pin)
* Node 326 = R8.2 (at pin)
* Node 264 = J10.7 (at pin)
* Node 327 = R7.2 (at pin)
* Node 270 = J10.6 (at pin)
* Node 328 = R6.2 (at pin)
* Node 276 = J10.5 (at pin)
* Node 329 = R5.2 (at pin)
* Node 282 = J10.4 (at pin)
* Node 330 = R4.2 (at pin)
* Node 288 = J10.3 (at pin)
* Node 331 = R3.2 (at pin)
* Node 294 = J10.2 (at pin)
* Node 332 = R2.2 (at pin)
* Node 296 = U1.AM10 (at pin) (driver)
X_mdl_297 297 Vinp MODEL_U1_AM10_ip
* Node 301 = J10.1 (at pin)

* Node   0 = Gnd (Common Return)

.connect 303 120 

.connect 319 216 

.connect 318 210 

.connect 317 204 

.connect 316 198 

.connect 315 192 

.connect 314 186 

.connect 313 180 

.connect 312 174 

.connect 311 168 

.connect 310 162 

.connect 309 156 

.connect 308 150 

.connect 307 144 

.connect 306 138 

.connect 305 132 

.connect 304 126 

.connect 332 294 

.connect 331 288 

.connect 330 282 

.connect 329 276 

.connect 328 270 

.connect 327 264 

.connect 326 258 

.connect 325 252 

.connect 324 246 

.connect 323 240 

.connect 322 234 

.connect 321 228 

.connect 320 222 


T001        101    0  106    0 Z0=5.983340e+001 TD=1.348640e-010
T002        101    0  104    0 Z0=5.000000e+001 TD=2.000000e-011
T003        101    0  105    0 Z0=5.000000e+001 TD=2.000000e-011
CP101       101    0 6.815e-014
REBD-J8_R102_2  106  108 22
TP102       104    0  109    0 Z0=1.092906e+002 TD=1.967232e-011
TP103       105    0  111    0 Z0=1.130906e+002 TD=2.148721e-011
T004        108    0  114    0 Z0=5.983340e+001 TD=2.252790e-011
R32_2       120    0 50
R31_2       126    0 50
R30_2       132    0 50
R29_2       138    0 50
R28_2       144    0 50
R27_2       150    0 50
R26_2       156    0 50
R25_2       162    0 50
R24_2       168    0 50
R23_2       174    0 50
R22_2       180    0 50
R21_2       186    0 50
R20_2       192    0 50
R19_2       198    0 50
R18_2       204    0 50
R16_2       210    0 50
R15_2       216    0 50
R14_2       222    0 50
R13_2       228    0 50
R12_2       234    0 50
R11_2       240    0 50
R10_2       246    0 50
R9_2        252    0 50
R8_2        258    0 50
R7_2        264    0 50
R6_2        270    0 50
R5_2        276    0 50
R4_2        282    0 50
R3_2        288    0 50
R2_2        294    0 50
TP195       296    0  297    0 Z0=1.013434e+002 TD=1.064105e-010
T005        296    0  299    0 Z0=4.333806e+001 TD=1.150930e-011
CV001       296    0 2.185e-014
W006       N=1  301    0  299    0 RLGCmodel=Model_W006 L=0.0972069 fgd=1e9  MULTIDEBYE=1
CV002       299    0 4.790e-013

V3  3  0  1.00
V2  2  0  1.80
V1  1  0  0.00

****  Transmission line models ***********************

*********************************
* Single uncoupled transmission line

.MODEL Model_W006 W MODELTYPE=RLGC N=1
* Lo  (H/m)
+ Lo =
+ 3.39994e-007

* Co  (F/m)
+ Co =
+ 1.30903e-010

* Ro (Ohm/m)
+ Ro =
+ 10.0819

* Go (S/m)
+ Go =
+ 0

* Rs (Ohm/m-sqrt(Hz))
+ Rs =
+ 0.00188059

* Gd (S/m-Hz)
+ Gd =
+ 1.64497e-011

****  End Transmission line models *******************

.ENDS

* IBIS model subcircuit definitions
**********************************************
*Define subcircuit for MODEL_EBD-J8_U15_J9_ip
.subckt MODEL_EBD-J8_U15_J9_ip a_signal d_receive 
VPullUpRef a_PURef 0 1.8
VPullDownRef a_PDRef 0 0

X_104 a_signal d_receive 0 a_PURef a_PDRef MODEL_EBD-J8_U15_J9

.ends MODEL_EBD-J8_U15_J9_ip

*Define subcircuit for MODEL_EBD-J8_U15_J9
.subckt MODEL_EBD-J8_U15_J9 a_signal d_receive a_gnd a_PURef a_PDRef 

C_comp a_signal a_gnd 2.811e-012

VGCRef a_GCRef 0 0
G_gnd_clamp a_signal a_GCRef table v(a_signal, a_GCRef) = 
+ (-23.4,-22.2654) (-1.8,-0.760219) (-1.795,-0.755241) 
+ (-1.79,-0.750299) (-1.785,-0.745359) (-1.78,-0.740421) 
+ (-1.775,-0.735484) (-1.77,-0.730549) (-1.765,-0.725617) 
+ (-1.755,-0.715754) (-1.735,-0.696055) (-1.73,-0.691139) 
+ (-1.695,-0.656751) (-1.69,-0.651848) (-1.63,-0.593191) 
+ (-1.625,-0.588303) (-1.62,-0.583444) (-1.615,-0.578597) 
+ (-1.55,-0.51558) (-1.545,-0.510732) (-1.54,-0.505913) 
+ (-1.53,-0.496355) (-1.525,-0.491576) (-1.45,-0.419894) 
+ (-1.445,-0.415115) (-1.44,-0.410336) (-1.435,-0.40558) 
+ (-1.415,-0.387037) (-1.41,-0.382402) (-1.32,-0.29896) 
+ (-1.315,-0.294325) (-1.3,-0.280418) (-1.295,-0.275794) 
+ (-1.27,-0.254226) (-1.265,-0.249912) (-1.175,-0.172264) 
+ (-1.17,-0.16795) (-1.16,-0.159323) (-1.155,-0.155515) 
+ (-1.14,-0.145365) (-1.135,-0.141982) (-1.04,-0.0776975) 
+ (-1.035,-0.0743141) (-1.01,-0.0573972) (-1.005,-0.0557414) 
+ (-0.98,-0.0484965) (-0.975,-0.0470476) (-0.94,-0.0369047) 
+ (-0.935,-0.0354557) (-0.895,-0.0238639) (-0.89,-0.0230547) 
+ (-0.875,-0.0215177) (-0.87,-0.0210053) (-0.825,-0.0163943) 
+ (-0.82,-0.0158819) (-0.795,-0.0133202) (-0.79,-0.0128917) 
+ (-0.78,-0.0122114) (-0.775,-0.0118712) (-0.745,-0.00983015) 
+ (-0.74,-0.00948997) (-0.7,-0.00676859) (-0.695,-0.0065163) 
+ (-0.69,-0.00628185) (-0.685,-0.0060474) (-0.65,-0.00440625) 
+ (-0.645,-0.00417181) (-0.615,-0.00276511) (-0.61,-0.00255864) 
+ (-0.605,-0.0024436) (-0.56,-0.00140824) (-0.555,-0.0012932) 
+ (-0.535,-0.000833048) (-0.53,-0.000718009) (-0.525,-0.00064001) 
+ (-0.515,-0.000581028) (-0.51,-0.000551537) (-0.49,-0.000433574) 
+ (-0.485,-0.000404083) (-0.475,-0.000345101) (-0.47,-0.00031561) 
+ (-0.44,-0.000138664) (-0.435,-0.000122592) (-0.41,-9.27216e-005) 
+ (-0.39,-6.88249e-005) (-0.385,-6.50985e-005) (-0.365,-5.80787e-005) 
+ (-0.355,-5.45688e-005) (-0.35,-5.28139e-005) (-0.325,-4.40391e-005) 
+ (-0.32,-4.25496e-005) (-0.285,0) (3.6,0) 
+ (25.2,0) 

VPCRef a_PCRef 0 1.8
G_power_clamp a_PCRef a_signal table v(a_PCRef, a_signal) = 
+ (-23.4,-18.3) (-1.8,-0.607667) (-1.795,-0.603572) 
+ (-1.79,-0.599504) (-1.785,-0.595438) (-1.78,-0.591374) 
+ (-1.775,-0.587311) (-1.77,-0.58325) (-1.765,-0.57919) 
+ (-1.755,-0.571074) (-1.735,-0.554862) (-1.73,-0.550816) 
+ (-1.695,-0.522518) (-1.69,-0.518485) (-1.63,-0.470223) 
+ (-1.625,-0.466201) (-1.62,-0.462204) (-1.615,-0.458217) 
+ (-1.55,-0.406381) (-1.545,-0.402394) (-1.54,-0.39843) 
+ (-1.53,-0.390572) (-1.525,-0.386643) (-1.45,-0.327709) 
+ (-1.445,-0.32378) (-1.44,-0.319851) (-1.435,-0.315941) 
+ (-1.415,-0.300718) (-1.41,-0.296913) (-1.32,-0.228411) 
+ (-1.315,-0.224606) (-1.3,-0.213189) (-1.295,-0.209394) 
+ (-1.27,-0.191808) (-1.265,-0.188291) (-1.175,-0.124981) 
+ (-1.17,-0.121464) (-1.16,-0.114429) (-1.155,-0.111406) 
+ (-1.14,-0.103581) (-1.135,-0.100972) (-1.04,-0.0514083) 
+ (-1.035,-0.0487997) (-1.01,-0.0357566) (-1.005,-0.0346027) 
+ (-0.98,-0.0297033) (-0.975,-0.0287235) (-0.94,-0.0218644) 
+ (-0.935,-0.0208845) (-0.895,-0.0130456) (-0.89,-0.0124844) 
+ (-0.875,-0.0113837) (-0.87,-0.0110168) (-0.825,-0.0077146) 
+ (-0.82,-0.0073477) (-0.795,-0.00551317) (-0.79,-0.00523633) 
+ (-0.78,-0.00487255) (-0.775,-0.00469066) (-0.745,-0.00359931) 
+ (-0.74,-0.00341742) (-0.7,-0.0019623) (-0.695,-0.00186186) 
+ (-0.69,-0.00177795) (-0.685,-0.00169404) (-0.65,-0.00110668) 
+ (-0.645,-0.00102277) (-0.615,-0.000519312) (-0.61,-0.000449671) 
+ (-0.605,-0.000426662) (-0.56,-0.000219585) (-0.555,-0.000196577) 
+ (-0.535,-0.000104543) (-0.53,-8.15342e-005) (-0.525,-6.69439e-005) 
+ (-0.515,-5.98123e-005) (-0.51,-5.62465e-005) (-0.49,-4.19832e-005) 
+ (-0.475,-3.12858e-005) (-0.47,-2.77199e-005) (-0.44,-6.32505e-006) 
+ (-0.435,-4.48769e-006) (-0.41,-1.80397e-006) (-0.393,0) 
+ (3.6,0) (25.2,0) 

* IBIS style receiver logic.  No hysteresis.
Y_rx_logic ibis_receiver_logic(icx_behavioral)
+ GENERIC: corner="ibis_typ"
+          vinL_values="(0.650000,0.650000,0.650000)"
+          vinH_values="(1.150000,1.150000,1.150000)"
+ PORT: a_gnd
+       a_signal
+       d_receive

.model ibis_receiver_logic(icx_behavioral) MACRO LANG=VHDLAMS LIB=icxbase
.ends MODEL_EBD-J8_U15_J9

*Define subcircuit for MODEL_EBD-J8_U5_J1_ip
.subckt MODEL_EBD-J8_U5_J1_ip a_signal d_receive 
VPullUpRef a_PURef 0 1.8
VPullDownRef a_PDRef 0 0

X_105 a_signal d_receive 0 a_PURef a_PDRef MODEL_EBD-J8_U5_J1

.ends MODEL_EBD-J8_U5_J1_ip

*Define subcircuit for MODEL_EBD-J8_U5_J1
.subckt MODEL_EBD-J8_U5_J1 a_signal d_receive a_gnd a_PURef a_PDRef 

C_comp a_signal a_gnd 2.811e-012

VGCRef a_GCRef 0 0
G_gnd_clamp a_signal a_GCRef table v(a_signal, a_GCRef) = 
+ (-23.4,-22.2654) (-1.8,-0.760219) (-1.795,-0.755241) 
+ (-1.79,-0.750299) (-1.785,-0.745359) (-1.78,-0.740421) 
+ (-1.775,-0.735484) (-1.77,-0.730549) (-1.765,-0.725617) 
+ (-1.755,-0.715754) (-1.735,-0.696055) (-1.73,-0.691139) 
+ (-1.695,-0.656751) (-1.69,-0.651848) (-1.63,-0.593191) 
+ (-1.625,-0.588303) (-1.62,-0.583444) (-1.615,-0.578597) 
+ (-1.55,-0.51558) (-1.545,-0.510732) (-1.54,-0.505913) 
+ (-1.53,-0.496355) (-1.525,-0.491576) (-1.45,-0.419894) 
+ (-1.445,-0.415115) (-1.44,-0.410336) (-1.435,-0.40558) 
+ (-1.415,-0.387037) (-1.41,-0.382402) (-1.32,-0.29896) 
+ (-1.315,-0.294325) (-1.3,-0.280418) (-1.295,-0.275794) 
+ (-1.27,-0.254226) (-1.265,-0.249912) (-1.175,-0.172264) 
+ (-1.17,-0.16795) (-1.16,-0.159323) (-1.155,-0.155515) 
+ (-1.14,-0.145365) (-1.135,-0.141982) (-1.04,-0.0776975) 
+ (-1.035,-0.0743141) (-1.01,-0.0573972) (-1.005,-0.0557414) 
+ (-0.98,-0.0484965) (-0.975,-0.0470476) (-0.94,-0.0369047) 
+ (-0.935,-0.0354557) (-0.895,-0.0238639) (-0.89,-0.0230547) 
+ (-0.875,-0.0215177) (-0.87,-0.0210053) (-0.825,-0.0163943) 
+ (-0.82,-0.0158819) (-0.795,-0.0133202) (-0.79,-0.0128917) 
+ (-0.78,-0.0122114) (-0.775,-0.0118712) (-0.745,-0.00983015) 
+ (-0.74,-0.00948997) (-0.7,-0.00676859) (-0.695,-0.0065163) 
+ (-0.69,-0.00628185) (-0.685,-0.0060474) (-0.65,-0.00440625) 
+ (-0.645,-0.00417181) (-0.615,-0.00276511) (-0.61,-0.00255864) 
+ (-0.605,-0.0024436) (-0.56,-0.00140824) (-0.555,-0.0012932) 
+ (-0.535,-0.000833048) (-0.53,-0.000718009) (-0.525,-0.00064001) 
+ (-0.515,-0.000581028) (-0.51,-0.000551537) (-0.49,-0.000433574) 
+ (-0.485,-0.000404083) (-0.475,-0.000345101) (-0.47,-0.00031561) 
+ (-0.44,-0.000138664) (-0.435,-0.000122592) (-0.41,-9.27216e-005) 
+ (-0.39,-6.88249e-005) (-0.385,-6.50985e-005) (-0.365,-5.80787e-005) 
+ (-0.355,-5.45688e-005) (-0.35,-5.28139e-005) (-0.325,-4.40391e-005) 
+ (-0.32,-4.25496e-005) (-0.285,0) (3.6,0) 
+ (25.2,0) 

VPCRef a_PCRef 0 1.8
G_power_clamp a_PCRef a_signal table v(a_PCRef, a_signal) = 
+ (-23.4,-18.3) (-1.8,-0.607667) (-1.795,-0.603572) 
+ (-1.79,-0.599504) (-1.785,-0.595438) (-1.78,-0.591374) 
+ (-1.775,-0.587311) (-1.77,-0.58325) (-1.765,-0.57919) 
+ (-1.755,-0.571074) (-1.735,-0.554862) (-1.73,-0.550816) 
+ (-1.695,-0.522518) (-1.69,-0.518485) (-1.63,-0.470223) 
+ (-1.625,-0.466201) (-1.62,-0.462204) (-1.615,-0.458217) 
+ (-1.55,-0.406381) (-1.545,-0.402394) (-1.54,-0.39843) 
+ (-1.53,-0.390572) (-1.525,-0.386643) (-1.45,-0.327709) 
+ (-1.445,-0.32378) (-1.44,-0.319851) (-1.435,-0.315941) 
+ (-1.415,-0.300718) (-1.41,-0.296913) (-1.32,-0.228411) 
+ (-1.315,-0.224606) (-1.3,-0.213189) (-1.295,-0.209394) 
+ (-1.27,-0.191808) (-1.265,-0.188291) (-1.175,-0.124981) 
+ (-1.17,-0.121464) (-1.16,-0.114429) (-1.155,-0.111406) 
+ (-1.14,-0.103581) (-1.135,-0.100972) (-1.04,-0.0514083) 
+ (-1.035,-0.0487997) (-1.01,-0.0357566) (-1.005,-0.0346027) 
+ (-0.98,-0.0297033) (-0.975,-0.0287235) (-0.94,-0.0218644) 
+ (-0.935,-0.0208845) (-0.895,-0.0130456) (-0.89,-0.0124844) 
+ (-0.875,-0.0113837) (-0.87,-0.0110168) (-0.825,-0.0077146) 
+ (-0.82,-0.0073477) (-0.795,-0.00551317) (-0.79,-0.00523633) 
+ (-0.78,-0.00487255) (-0.775,-0.00469066) (-0.745,-0.00359931) 
+ (-0.74,-0.00341742) (-0.7,-0.0019623) (-0.695,-0.00186186) 
+ (-0.69,-0.00177795) (-0.685,-0.00169404) (-0.65,-0.00110668) 
+ (-0.645,-0.00102277) (-0.615,-0.000519312) (-0.61,-0.000449671) 
+ (-0.605,-0.000426662) (-0.56,-0.000219585) (-0.555,-0.000196577) 
+ (-0.535,-0.000104543) (-0.53,-8.15342e-005) (-0.525,-6.69439e-005) 
+ (-0.515,-5.98123e-005) (-0.51,-5.62465e-005) (-0.49,-4.19832e-005) 
+ (-0.475,-3.12858e-005) (-0.47,-2.77199e-005) (-0.44,-6.32505e-006) 
+ (-0.435,-4.48769e-006) (-0.41,-1.80397e-006) (-0.393,0) 
+ (3.6,0) (25.2,0) 

* IBIS style receiver logic.  No hysteresis.
Y_rx_logic ibis_receiver_logic(icx_behavioral)
+ GENERIC: corner="ibis_typ"
+          vinL_values="(0.650000,0.650000,0.650000)"
+          vinH_values="(1.150000,1.150000,1.150000)"
+ PORT: a_gnd
+       a_signal
+       d_receive

.model ibis_receiver_logic(icx_behavioral) MACRO LANG=VHDLAMS LIB=icxbase
.ends MODEL_EBD-J8_U5_J1

*Define subcircuit for MODEL_U1_AM10_ip
.subckt MODEL_U1_AM10_ip a_signal a_control 
VPullUpRef a_PURef 0 1.8
VPullDownRef a_PDRef 0 1e-100


Y_a_control ibis_driver_logic(icx_behavioral)
+ GENERIC: corner="ibis_typ"
+          vmeas_values="( 0.5, 0.5, 0.5 )"
+ PORT: a_control
+       a_gnd
+       d_control

.model ibis_driver_logic(icx_behavioral) MACRO LANG=VHDLAMS LIB=icxbase

X_296 a_signal d_control 0 a_PURef a_PDRef MODEL_U1_AM10

.ends MODEL_U1_AM10_ip

*Define subcircuit for MODEL_U1_AM10
.subckt MODEL_U1_AM10 a_signal d_control a_gnd a_PURef a_PDRef

C_comp a_signal a_gnd 2.29e-012

VGCRef a_GCRef 0 0
G_gnd_clamp a_signal a_GCRef table v(a_signal, a_GCRef) = 
+ (-16.2,-531.037) (-1.8,-38.881) (-1.76,-37.5139) 
+ (-1.72,-36.1404) (-1.68,-35.37) (-1.64,-34.48) 
+ (-1.6,-33.864) (-1.56,-32.7827) (-1.52,-31.213) 
+ (-1.48,-30.43) (-1.44,-29.96) (-1.4,-28.362) 
+ (-1.36,-27.192) (-1.32,-26.326) (-1.28,-25.27) 
+ (-1.24,-24.56) (-1.2,-6.859) (-1.16,-1.998) 
+ (-1.12,-0.6476) (-1.08,-0.2564) (-1.04,-0.1286) 
+ (-1,-0.07477) (-0.96,-0.04437) (-0.92,-0.02541) 
+ (-0.88,-0.01527) (-0.84,-0.01068) (-0.8,-0.00833) 
+ (-0.76,-0.006779) (-0.72,-0.005583) (-0.68,-0.00455) 
+ (-0.64,-0.003606) (-0.6,-0.00274) (-0.56,-0.001965) 
+ (-0.52,-0.001303) (-0.48,-0.0007803) (-0.44,-0.0004131) 
+ (-0.4,-0.0001921) (-0.36,-7.91e-005) (-0.32,-2.898e-005) 
+ (-0.28,-9.395e-006) (-0.24,-2.701e-006) (-0.2,-7.023e-007) 
+ (-0.16,-1.693e-007) (-0.12,-3.87e-008) (-0.08,-8.68e-009) 
+ (-0.04,-8.505e-009) (0.24,-3.814e-010) (0.28,-1.765e-010) 
+ (0.32,-1.331e-010) (0.36,-9.055e-011) (0.4,-4.862e-011) 
+ (0.44,-7.086e-012) (0.48,3.416e-011) (0.52,7.522e-011) 
+ (0.56,1.161e-010) (0.6,1.57e-010) (0.64,1.977e-010) 
+ (0.68,2.384e-010) (0.72,2.791e-010) (0.76,3.198e-010) 
+ (0.8,3.605e-010) (0.84,4.013e-010) (0.88,4.421e-010) 
+ (0.92,4.83e-010) (0.96,5.239e-010) (1,5.649e-010) 
+ (1.04,6.06e-010) (1.08,6.472e-010) (1.12,6.886e-010) 
+ (1.16,7.301e-010) (1.2,7.717e-010) (1.24,8.135e-010) 
+ (1.28,8.555e-010) (1.32,8.977e-010) (1.36,9.402e-010) 
+ (1.4,9.83e-010) (1.44,1.026e-009) (1.48,1.069e-009) 
+ (1.52,1.11e-009) (1.56,1.148e-009) (1.6,1.181e-009) 
+ (1.64,1.214e-009) (1.68,1.25e-009) (1.72,1.3e-009) 
+ (1.76,1.389e-009) (1.8,1.595e-009) (16.2,7.5755e-008) 

VPCRef a_PCRef 0 1.8
G_power_clamp a_PCRef a_signal table v(a_PCRef, a_signal) = 
+ (-9,-5.892) (-1.8,-0.636) (-1.78,-0.6214) 
+ (-1.76,-0.6068) (-1.74,-0.5922) (-1.72,-0.5775) 
+ (-1.7,-0.5629) (-1.68,-0.5483) (-1.66,-0.5337) 
+ (-1.64,-0.5191) (-1.62,-0.5045) (-1.6,-0.4899) 
+ (-1.58,-0.4753) (-1.56,-0.4608) (-1.54,-0.4462) 
+ (-1.52,-0.4317) (-1.5,-0.4173) (-1.48,-0.4029) 
+ (-1.46,-0.3885) (-1.44,-0.3741) (-1.42,-0.3598) 
+ (-1.4,-0.3455) (-1.38,-0.3312) (-1.36,-0.3169) 
+ (-1.34,-0.3026) (-1.32,-0.2884) (-1.3,-0.2741) 
+ (-1.28,-0.2599) (-1.26,-0.2458) (-1.24,-0.2317) 
+ (-1.22,-0.2176) (-1.2,-0.2035) (-1.18,-0.1895) 
+ (-1.16,-0.1755) (-1.14,-0.1616) (-1.12,-0.1478) 
+ (-1.1,-0.1341) (-1.08,-0.1205) (-1.06,-0.107) 
+ (-1.04,-0.09377) (-1.02,-0.08082) (-1,-0.06827) 
+ (-0.98,-0.05627) (-0.96,-0.04504) (-0.94,-0.03489) 
+ (-0.92,-0.02617) (-0.9,-0.01921) (-0.88,-0.01418) 
+ (-0.86,-0.01087) (-0.84,-0.008828) (-0.82,-0.007559) 
+ (-0.8,-0.006709) (-0.78,-0.00607) (-0.76,-0.005538) 
+ (-0.74,-0.00506) (-0.72,-0.004614) (-0.7,-0.004188) 
+ (-0.68,-0.003778) (-0.66,-0.003383) (-0.64,-0.003003) 
+ (-0.62,-0.002638) (-0.6,-0.00229) (-0.58,-0.00196) 
+ (-0.56,-0.00165) (-0.54,-0.001363) (-0.52,-0.001101) 
+ (-0.5,-0.0008655) (-0.48,-0.00066) (-0.46,-0.000486) 
+ (-0.44,-0.0003443) (-0.42,-0.000234) (-0.4,-0.0001527) 
+ (-0.38,-9.58e-005) (-0.36,-5.812e-005) (-0.34,-3.427e-005) 
+ (-0.32,-1.972e-005) (-0.3,-1.11e-005) (-0.28,-6.116e-006) 
+ (-0.26,-3.299e-006) (-0.24,-1.743e-006) (-0.22,-9.032e-007) 
+ (-0.2,-4.598e-007) (-0.18,-2.305e-007) (-0.16,-1.14e-007) 
+ (-0.14,-5.589e-008) (-0.12,-2.735e-008) (-0.1,-1.354e-008) 
+ (-0.08,-6.966e-009) (-0.06,-3.891e-009) (-0.04,-2.482e-009) 
+ (-0.02,-1.857e-009) (0,-1.595e-009) (7.2,9.2725e-008) 

Y_control ibis_control(icx_behavioral)
+ PORT: d_control
+       d_pullup_control
+       d_pulldown_control

.model ibis_control(icx_behavioral) MACRO LANG=VHDLAMS LIB=icxbase


*IBIS Pulldown tables
Y_PullDown ibis_ktiv(icx_behavioral)
+ GENERIC: corner="ibis_typ"
+          tdata_0to1_typ="(4.96516e-012, 1.23871e-011, 1.9809e-011, 2.7231e-011, 3.46529e-011, 4.20748e-011,
+ 4.94968e-011, 5.69187e-011, 6.43406e-011, 7.17626e-011, 7.91845e-011, 8.66065e-011,
+ 9.40284e-011, 1.0145e-010, 1.08872e-010, 1.16294e-010, 1.23716e-010, 1.31138e-010,
+ 1.3856e-010, 1.45982e-010, 1.53404e-010, 1.60826e-010, 1.68248e-010, 1.7567e-010,
+ 1.83092e-010, 1.90514e-010, 1.97935e-010, 2.05357e-010, 2.12779e-010, 2.20201e-010,
+ 2.27623e-010, 2.35045e-010, 2.42467e-010, 2.49889e-010, 2.57311e-010, 2.64733e-010,
+ 2.72155e-010, 2.79577e-010, 2.86999e-010, 2.94421e-010, 3.01843e-010, 3.09265e-010,
+ 3.16686e-010, 3.24108e-010, 3.3153e-010, 3.38952e-010, 3.46374e-010, 3.53796e-010,
+ 3.61218e-010, 3.6864e-010, 3.76062e-010, 3.83484e-010, 3.90906e-010, 3.98328e-010,
+ 4.0575e-010, 4.13172e-010, 4.20594e-010, 4.28015e-010, 4.35437e-010, 4.42859e-010,
+ 4.50281e-010, 4.57703e-010, 4.65125e-010, 4.72547e-010, 4.79969e-010, 4.87391e-010,
+ 4.94813e-010, 5.02235e-010, 5.09657e-010, 5.17079e-010, 5.24501e-010, 5.31923e-010,
+ 5.39345e-010, 5.46766e-010, 5.54188e-010, 5.6161e-010, 5.69032e-010, 5.76454e-010,
+ 5.83876e-010, 5.91298e-010, 5.9872e-010, 6.06142e-010, 6.13564e-010, 6.20986e-010,
+ 6.28408e-010, 6.3583e-010, 6.43252e-010, 6.50674e-010, 6.58095e-010, 6.65517e-010,
+ 6.72939e-010, 6.80361e-010, 6.87783e-010, 6.95205e-010, 7.02627e-010, 7.10049e-010,
+ 7.17471e-010, 7.24893e-010, 7.32315e-010, 7.39737e-010, 7.47159e-010, 7.54581e-010,
+ 7.62003e-010, 7.69425e-010, 7.76846e-010, 7.84268e-010, 7.9169e-010, 7.99112e-010,
+ 8.06534e-010, 8.13956e-010, 8.21378e-010, 8.288e-010, 8.36222e-010, 8.43644e-010,
+ 8.51066e-010, 8.58488e-010, 8.6591e-010, 8.73332e-010, 8.80754e-010, 8.88175e-010,
+ 8.95597e-010, 9.03019e-010, 9.10441e-010, 9.17863e-010, 9.25285e-010, 9.32707e-010,
+ 9.40129e-010, 9.47551e-010, 9.54973e-010, 9.62395e-010, 9.69817e-010, 9.77239e-010,
+ 9.84661e-010, 9.92083e-010, 9.99505e-010, 1.00693e-009, 1.01435e-009, 1.02177e-009,
+ 1.02919e-009, 1.03661e-009, 1.04404e-009, 1.05146e-009, 1.05888e-009, 1.0663e-009,
+ 1.07372e-009, 1.08115e-009, 1.08857e-009, 1.09599e-009, 1.10341e-009, 1.11083e-009,
+ 1.11826e-009, 1.12568e-009, 1.1331e-009, 1.14052e-009, 1.14794e-009, 1.15537e-009,
+ 1.16279e-009, 1.17021e-009, 1.17763e-009, 1.18505e-009, 1.19247e-009, 1.1999e-009,
+ 1.20732e-009, 1.21474e-009, 1.22216e-009, 1.22958e-009, 1.23701e-009, 1.24443e-009,
+ 1.25185e-009, 1.25927e-009, 1.26669e-009, 1.27412e-009, 1.28154e-009, 1.28896e-009,
+ 1.29638e-009, 1.3038e-009, 1.31123e-009, 1.31865e-009, 1.32607e-009, 1.33349e-009,
+ 1.34091e-009, 1.34834e-009, 1.35576e-009, 1.36318e-009, 1.3706e-009, 1.37802e-009,
+ 1.38545e-009, 1.39287e-009, 1.40029e-009, 1.40771e-009, 1.41513e-009, 1.42255e-009,
+ 1.42998e-009, 1.4374e-009, 1.44482e-009, 1.45224e-009, 1.45966e-009, 1.46709e-009,
+ 1.47451e-009, 1.48193e-009, 1.48935e-009, 1.49677e-009, 1.5042e-009)"
+          kdata_0to1_typ="(0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0.00569651, 0.00797394, 0.0101697, 0.0122872, 0.0456626,
+ 0.0510044, 0.0561412, 0.0610819, 0.0899824, 0.0974826, 0.104784,
+ 0.111894, 0.118823, 0.177096, 0.188923, 0.200394, 0.211537,
+ 0.222298, 0.255786, 0.267891, 0.279519, 0.290826, 0.345133,
+ 0.360612, 0.375734, 0.390569, 0.424544, 0.441794, 0.458924,
+ 0.475911, 0.515607, 0.53587, 0.556206, 0.576611, 0.596363,
+ 0.618281, 0.640704, 0.663382, 0.663809, 0.684793, 0.706227,
+ 0.728215, 0.739928, 0.762191, 0.784981, 0.808267, 0.781378,
+ 0.798831, 0.816575, 0.834617, 0.837009, 0.853991, 0.871298,
+ 0.888938, 0.853994, 0.864319, 0.87483, 0.885447, 0.896391,
+ 0.907642, 0.919051, 0.930624, 0.915004, 0.922767, 0.930609,
+ 0.93853, 0.935223, 0.941614, 0.948057, 0.954555, 0.943771,
+ 0.947669, 0.951587, 0.955524, 0.954325, 0.957495, 0.960677,
+ 0.963872, 0.959697, 0.961761, 0.96383, 0.965904, 0.965428,
+ 0.96711, 0.968795, 0.970484, 0.969038, 0.970237, 0.971437,
+ 0.97264, 0.973112, 0.974201, 0.975292, 0.976383, 0.975782,
+ 0.976605, 0.977428, 0.978253, 0.980456, 0.981505, 0.982555,
+ 0.983607, 0.982997, 0.98378, 0.984564, 0.985349, 0.984822,
+ 0.985393, 0.985964, 0.986536, 0.986131, 0.986543, 0.986954,
+ 0.987366, 0.987778, 0.987452, 0.987759, 0.988067, 0.988374,
+ 0.988708, 0.989019, 0.989331, 0.989643, 0.989984, 0.990301,
+ 0.990617, 0.990934, 0.990885, 0.991149, 0.991413, 0.991677,
+ 0.991961, 0.992228, 0.992495, 0.992763, 0.992662, 0.992875,
+ 0.993089, 0.993302, 0.994259, 0.994583, 0.994907, 0.995231,
+ 0.994741, 0.994944, 0.995147, 0.99535, 0.995553, 0.995502,
+ 0.995665, 0.995828, 0.995991, 0.995808, 0.995915, 0.996023,
+ 0.996131, 0.996242, 0.99635, 0.996458, 0.996566, 0.996678,
+ 0.996787, 0.996896, 0.997005, 0.997116, 0.997225, 0.997334,
+ 0.997444, 0.997555, 0.997665, 0.997775, 0.997885, 0.997657,
+ 0.997711, 0.997765, 0.997819, 0.997872, 1)"
+          tdata_1to0_typ="(2.10524e-010, 2.16774e-010, 2.23024e-010, 2.29274e-010, 2.35524e-010, 2.41774e-010,
+ 2.48024e-010, 2.54274e-010, 2.60524e-010, 2.66774e-010, 2.73024e-010, 2.79274e-010,
+ 2.85524e-010, 2.91774e-010, 2.98024e-010, 3.04274e-010, 3.10524e-010, 3.16774e-010,
+ 3.23024e-010, 3.29274e-010, 3.35524e-010, 3.41774e-010, 3.48024e-010, 3.54274e-010,
+ 3.60524e-010, 3.66774e-010, 3.73024e-010, 3.79274e-010, 3.85524e-010, 3.91774e-010,
+ 3.98024e-010, 4.04274e-010, 4.10524e-010, 4.16774e-010, 4.23024e-010, 4.29274e-010,
+ 4.35524e-010, 4.41774e-010, 4.48024e-010, 4.54274e-010, 4.60524e-010, 4.66774e-010,
+ 4.73024e-010, 4.79274e-010, 4.85524e-010, 4.91774e-010, 4.98024e-010, 5.04274e-010,
+ 5.10524e-010, 5.16774e-010, 5.23024e-010, 5.29274e-010, 5.35524e-010, 5.41774e-010,
+ 5.48024e-010, 5.54274e-010, 5.60524e-010, 5.66774e-010, 5.73024e-010, 5.79274e-010,
+ 5.85524e-010, 5.91774e-010, 5.98024e-010, 6.04274e-010, 6.10524e-010, 6.16774e-010,
+ 6.23024e-010, 6.29274e-010, 6.35524e-010, 6.41774e-010, 6.48024e-010, 6.54274e-010,
+ 6.60524e-010, 6.66774e-010, 6.73024e-010, 6.79274e-010, 6.85524e-010, 6.91774e-010,
+ 6.98024e-010, 7.04274e-010, 7.10524e-010, 7.16774e-010, 7.23024e-010, 7.29274e-010,
+ 7.35524e-010, 7.41774e-010, 7.48024e-010, 7.54274e-010, 7.60524e-010, 7.66774e-010,
+ 7.73024e-010, 7.79274e-010, 7.85524e-010, 7.91774e-010, 7.98024e-010, 8.04274e-010,
+ 8.10524e-010, 8.16774e-010, 8.23024e-010, 8.29274e-010, 8.35524e-010, 8.41774e-010,
+ 8.48024e-010, 8.54274e-010, 8.60524e-010, 8.66774e-010, 8.73024e-010, 8.79274e-010,
+ 8.85524e-010, 8.91774e-010, 8.98024e-010, 9.04274e-010, 9.10524e-010, 9.16774e-010,
+ 9.23024e-010, 9.29274e-010, 9.35524e-010, 9.41774e-010, 9.48024e-010, 9.54274e-010,
+ 9.60524e-010, 9.66774e-010, 9.73024e-010, 9.79274e-010, 9.85524e-010, 9.91774e-010,
+ 9.98024e-010, 1.00427e-009, 1.01052e-009, 1.01677e-009, 1.02302e-009, 1.02927e-009,
+ 1.03552e-009, 1.04177e-009, 1.04802e-009, 1.05427e-009, 1.06052e-009, 1.06677e-009,
+ 1.07302e-009, 1.07927e-009, 1.08552e-009, 1.09177e-009, 1.09802e-009, 1.10427e-009,
+ 1.11052e-009, 1.11677e-009, 1.12302e-009, 1.12927e-009, 1.13552e-009, 1.14177e-009,
+ 1.14802e-009, 1.15427e-009, 1.16052e-009, 1.16677e-009, 1.17302e-009, 1.17927e-009,
+ 1.18552e-009, 1.19177e-009, 1.19802e-009, 1.20427e-009, 1.21052e-009, 1.21677e-009,
+ 1.22302e-009, 1.22927e-009, 1.23552e-009, 1.24177e-009, 1.24802e-009, 1.25427e-009,
+ 1.26052e-009, 1.26677e-009, 1.27302e-009, 1.27927e-009, 1.28552e-009, 1.29177e-009,
+ 1.29802e-009, 1.30427e-009, 1.31052e-009, 1.31677e-009, 1.32302e-009, 1.32927e-009,
+ 1.33552e-009, 1.34177e-009, 1.34802e-009, 1.35427e-009, 1.36052e-009, 1.36677e-009,
+ 1.37302e-009, 1.37927e-009, 1.38552e-009, 1.39177e-009, 1.39802e-009, 1.40427e-009,
+ 1.41052e-009, 1.41677e-009, 1.42302e-009, 1.42927e-009, 1.43552e-009, 1.44177e-009,
+ 1.44802e-009, 1.45427e-009, 1.46052e-009, 1.46677e-009)"
+          kdata_1to0_typ="(1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 0.994646, 0.993826, 0.993007, 0.992189, 0.980394,
+ 0.978163, 0.975939, 0.973721, 0.97151, 0.945079, 0.939915,
+ 0.93477, 0.929645, 0.924539, 0.91305, 0.907394, 0.901718,
+ 0.896024, 0.890313, 0.817187, 0.80378, 0.790449, 0.777194,
+ 0.764017, 0.726053, 0.710242, 0.694453, 0.67869, 0.55545,
+ 0.528887, 0.502923, 0.477672, 0.452928, 0.441447, 0.417835,
+ 0.394483, 0.371407, 0.348571, 0.281799, 0.255858, 0.230407,
+ 0.20539, 0.180756, 0.195081, 0.173155, 0.151292, 0.129533,
+ 0.107868, 0.118215, 0.0991421, 0.0800503, 0.0609434, 0.0418339,
+ 0.0555166, 0.0392241, 0.0228697, 0.00641968, 0.0495123, 0.0386718,
+ 0.027634, 0.0164357, 0.00508082, 0.0142965, 0.00525532, 0,
+ 0, 0, 0.011854, 0.00700832, 0.00205821, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 5.24679e-005, 0.00025246,
+ 0.000453967, 0.000657004, 0.000861589, 0.00106774, 0.00127547, 0.0014848,
+ 0.00169204, 0.0019002, 0.00210928, 0.00231928, 0.00100161, 0.00100357,
+ 0.00100553, 0.0010075, 0.00100947, 0.00100465, 0.00100577, 0.00100691,
+ 0.00100804, 0.00100918, 0.00101032, 0.00101146, 0.0010126, 0.00101375,
+ 0.00101491, 0.00101366, 0.00101452, 0.00101539, 0.00101627, 0.00101714,
+ 0.00101553, 0.00101612, 0.0010167, 0.00101728, 0.00101787, 0.00101845,
+ 0.00101904, 0.00101962, 0.00102021, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0)"
+          vdata_typ="(-0.9, -0.84, -0.78, -0.72, -0.66, -0.6,
+ -0.54, -0.48, -0.42, -0.36, -0.3, -0.24,
+ -0.18, -0.12, -0.06, 0, 0.06, 0.12,
+ 0.18, 0.24, 0.3, 0.36, 0.42, 0.48,
+ 0.54, 0.6, 0.66, 0.72, 0.78, 0.84,
+ 0.9, 0.96, 1.02, 1.08, 1.14, 1.2,
+ 1.26, 1.32, 1.38, 1.44, 1.5, 1.56,
+ 1.62, 1.68, 1.74, 1.8, 1.86, 1.92,
+ 1.98, 2.04, 2.1, 2.16, 2.22, 2.28,
+ 2.34, 2.4, 2.46, 2.52, 2.58, 2.64,
+ 2.7, 2.76, 2.82, 2.88, 2.94, 3,
+ 3.06, 3.12, 3.18, 3.24, 3.3, 3.36,
+ 3.42, 3.48, 3.54, 3.6)"
+          idata_typ="(-0.02224, -0.02215, -0.021557, -0.020807, -0.019932, -0.01894,
+ -0.017762, -0.0163597, -0.0146538, -0.0127109, -0.0106332, -0.0085203,
+ -0.0063937, -0.004263, -0.002132, 0, 0.002124, 0.004233,
+ 0.006324, 0.008397, 0.01045, 0.01249, 0.0145, 0.01649,
+ 0.01846, 0.0204, 0.02231, 0.0242, 0.02606, 0.0279,
+ 0.0297, 0.03146, 0.0332, 0.03489, 0.03655, 0.03817,
+ 0.03974, 0.04128, 0.04276, 0.04419, 0.04556, 0.04688,
+ 0.04813, 0.04932, 0.05042, 0.05145, 0.05239, 0.05324,
+ 0.0539998, 0.0546683, 0.0552489, 0.0557519, 0.056186, 0.05657,
+ 0.056897, 0.0572, 0.057457, 0.057706, 0.05793, 0.058132,
+ 0.05833, 0.05856, 0.05869, 0.0588, 0.0591, 0.0592,
+ 0.0593, 0.0594, 0.0596, 0.0598, 0.0599, 0.06,
+ 0.0602, 0.0603, 0.0604, 0.0606)"
+          tdata_0to1_min="(4.96516e-012, 1.23871e-011, 1.9809e-011, 2.7231e-011, 3.46529e-011, 4.20748e-011,
+ 4.94968e-011, 5.69187e-011, 6.43406e-011, 7.17626e-011, 7.91845e-011, 8.66065e-011,
+ 9.40284e-011, 1.0145e-010, 1.08872e-010, 1.16294e-010, 1.23716e-010, 1.31138e-010,
+ 1.3856e-010, 1.45982e-010, 1.53404e-010, 1.60826e-010, 1.68248e-010, 1.7567e-010,
+ 1.83092e-010, 1.90514e-010, 1.97935e-010, 2.05357e-010, 2.12779e-010, 2.20201e-010,
+ 2.27623e-010, 2.35045e-010, 2.42467e-010, 2.49889e-010, 2.57311e-010, 2.64733e-010,
+ 2.72155e-010, 2.79577e-010, 2.86999e-010, 2.94421e-010, 3.01843e-010, 3.09265e-010,
+ 3.16686e-010, 3.24108e-010, 3.3153e-010, 3.38952e-010, 3.46374e-010, 3.53796e-010,
+ 3.61218e-010, 3.6864e-010, 3.76062e-010, 3.83484e-010, 3.90906e-010, 3.98328e-010,
+ 4.0575e-010, 4.13172e-010, 4.20594e-010, 4.28015e-010, 4.35437e-010, 4.42859e-010,
+ 4.50281e-010, 4.57703e-010, 4.65125e-010, 4.72547e-010, 4.79969e-010, 4.87391e-010,
+ 4.94813e-010, 5.02235e-010, 5.09657e-010, 5.17079e-010, 5.24501e-010, 5.31923e-010,
+ 5.39345e-010, 5.46766e-010, 5.54188e-010, 5.6161e-010, 5.69032e-010, 5.76454e-010,
+ 5.83876e-010, 5.91298e-010, 5.9872e-010, 6.06142e-010, 6.13564e-010, 6.20986e-010,
+ 6.28408e-010, 6.3583e-010, 6.43252e-010, 6.50674e-010, 6.58095e-010, 6.65517e-010,
+ 6.72939e-010, 6.80361e-010, 6.87783e-010, 6.95205e-010, 7.02627e-010, 7.10049e-010,
+ 7.17471e-010, 7.24893e-010, 7.32315e-010, 7.39737e-010, 7.47159e-010, 7.54581e-010,
+ 7.62003e-010, 7.69425e-010, 7.76846e-010, 7.84268e-010, 7.9169e-010, 7.99112e-010,
+ 8.06534e-010, 8.13956e-010, 8.21378e-010, 8.288e-010, 8.36222e-010, 8.43644e-010,
+ 8.51066e-010, 8.58488e-010, 8.6591e-010, 8.73332e-010, 8.80754e-010, 8.88175e-010,
+ 8.95597e-010, 9.03019e-010, 9.10441e-010, 9.17863e-010, 9.25285e-010, 9.32707e-010,
+ 9.40129e-010, 9.47551e-010, 9.54973e-010, 9.62395e-010, 9.69817e-010, 9.77239e-010,
+ 9.84661e-010, 9.92083e-010, 9.99505e-010, 1.00693e-009, 1.01435e-009, 1.02177e-009,
+ 1.02919e-009, 1.03661e-009, 1.04404e-009, 1.05146e-009, 1.05888e-009, 1.0663e-009,
+ 1.07372e-009, 1.08115e-009, 1.08857e-009, 1.09599e-009, 1.10341e-009, 1.11083e-009,
+ 1.11826e-009, 1.12568e-009, 1.1331e-009, 1.14052e-009, 1.14794e-009, 1.15537e-009,
+ 1.16279e-009, 1.17021e-009, 1.17763e-009, 1.18505e-009, 1.19247e-009, 1.1999e-009,
+ 1.20732e-009, 1.21474e-009, 1.22216e-009, 1.22958e-009, 1.23701e-009, 1.24443e-009,
+ 1.25185e-009, 1.25927e-009, 1.26669e-009, 1.27412e-009, 1.28154e-009, 1.28896e-009,
+ 1.29638e-009, 1.3038e-009, 1.31123e-009, 1.31865e-009, 1.32607e-009, 1.33349e-009,
+ 1.34091e-009, 1.34834e-009, 1.35576e-009, 1.36318e-009, 1.3706e-009, 1.37802e-009,
+ 1.38545e-009, 1.39287e-009, 1.40029e-009, 1.40771e-009, 1.41513e-009, 1.42255e-009,
+ 1.42998e-009, 1.4374e-009, 1.44482e-009, 1.45224e-009, 1.45966e-009, 1.46709e-009,
+ 1.47451e-009, 1.48193e-009, 1.48935e-009, 1.49677e-009, 1.5042e-009)"
+          kdata_0to1_min="(0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0.00569651, 0.00797394, 0.0101697, 0.0122872, 0.0456626,
+ 0.0510044, 0.0561412, 0.0610819, 0.0899824, 0.0974826, 0.104784,
+ 0.111894, 0.118823, 0.177096, 0.188923, 0.200394, 0.211537,
+ 0.222298, 0.255786, 0.267891, 0.279519, 0.290826, 0.345133,
+ 0.360612, 0.375734, 0.390569, 0.424544, 0.441794, 0.458924,
+ 0.475911, 0.515607, 0.53587, 0.556206, 0.576611, 0.596363,
+ 0.618281, 0.640704, 0.663382, 0.663809, 0.684793, 0.706227,
+ 0.728215, 0.739928, 0.762191, 0.784981, 0.808267, 0.781378,
+ 0.798831, 0.816575, 0.834617, 0.837009, 0.853991, 0.871298,
+ 0.888938, 0.853994, 0.864319, 0.87483, 0.885447, 0.896391,
+ 0.907642, 0.919051, 0.930624, 0.915004, 0.922767, 0.930609,
+ 0.93853, 0.935223, 0.941614, 0.948057, 0.954555, 0.943771,
+ 0.947669, 0.951587, 0.955524, 0.954325, 0.957495, 0.960677,
+ 0.963872, 0.959697, 0.961761, 0.96383, 0.965904, 0.965428,
+ 0.96711, 0.968795, 0.970484, 0.969038, 0.970237, 0.971437,
+ 0.97264, 0.973112, 0.974201, 0.975292, 0.976383, 0.975782,
+ 0.976605, 0.977428, 0.978253, 0.980456, 0.981505, 0.982555,
+ 0.983607, 0.982997, 0.98378, 0.984564, 0.985349, 0.984822,
+ 0.985393, 0.985964, 0.986536, 0.986131, 0.986543, 0.986954,
+ 0.987366, 0.987778, 0.987452, 0.987759, 0.988067, 0.988374,
+ 0.988708, 0.989019, 0.989331, 0.989643, 0.989984, 0.990301,
+ 0.990617, 0.990934, 0.990885, 0.991149, 0.991413, 0.991677,
+ 0.991961, 0.992228, 0.992495, 0.992763, 0.992662, 0.992875,
+ 0.993089, 0.993302, 0.994259, 0.994583, 0.994907, 0.995231,
+ 0.994741, 0.994944, 0.995147, 0.99535, 0.995553, 0.995502,
+ 0.995665, 0.995828, 0.995991, 0.995808, 0.995915, 0.996023,
+ 0.996131, 0.996242, 0.99635, 0.996458, 0.996566, 0.996678,
+ 0.996787, 0.996896, 0.997005, 0.997116, 0.997225, 0.997334,
+ 0.997444, 0.997555, 0.997665, 0.997775, 0.997885, 0.997657,
+ 0.997711, 0.997765, 0.997819, 0.997872, 1)"
+          tdata_1to0_min="(2.10524e-010, 2.16774e-010, 2.23024e-010, 2.29274e-010, 2.35524e-010, 2.41774e-010,
+ 2.48024e-010, 2.54274e-010, 2.60524e-010, 2.66774e-010, 2.73024e-010, 2.79274e-010,
+ 2.85524e-010, 2.91774e-010, 2.98024e-010, 3.04274e-010, 3.10524e-010, 3.16774e-010,
+ 3.23024e-010, 3.29274e-010, 3.35524e-010, 3.41774e-010, 3.48024e-010, 3.54274e-010,
+ 3.60524e-010, 3.66774e-010, 3.73024e-010, 3.79274e-010, 3.85524e-010, 3.91774e-010,
+ 3.98024e-010, 4.04274e-010, 4.10524e-010, 4.16774e-010, 4.23024e-010, 4.29274e-010,
+ 4.35524e-010, 4.41774e-010, 4.48024e-010, 4.54274e-010, 4.60524e-010, 4.66774e-010,
+ 4.73024e-010, 4.79274e-010, 4.85524e-010, 4.91774e-010, 4.98024e-010, 5.04274e-010,
+ 5.10524e-010, 5.16774e-010, 5.23024e-010, 5.29274e-010, 5.35524e-010, 5.41774e-010,
+ 5.48024e-010, 5.54274e-010, 5.60524e-010, 5.66774e-010, 5.73024e-010, 5.79274e-010,
+ 5.85524e-010, 5.91774e-010, 5.98024e-010, 6.04274e-010, 6.10524e-010, 6.16774e-010,
+ 6.23024e-010, 6.29274e-010, 6.35524e-010, 6.41774e-010, 6.48024e-010, 6.54274e-010,
+ 6.60524e-010, 6.66774e-010, 6.73024e-010, 6.79274e-010, 6.85524e-010, 6.91774e-010,
+ 6.98024e-010, 7.04274e-010, 7.10524e-010, 7.16774e-010, 7.23024e-010, 7.29274e-010,
+ 7.35524e-010, 7.41774e-010, 7.48024e-010, 7.54274e-010, 7.60524e-010, 7.66774e-010,
+ 7.73024e-010, 7.79274e-010, 7.85524e-010, 7.91774e-010, 7.98024e-010, 8.04274e-010,
+ 8.10524e-010, 8.16774e-010, 8.23024e-010, 8.29274e-010, 8.35524e-010, 8.41774e-010,
+ 8.48024e-010, 8.54274e-010, 8.60524e-010, 8.66774e-010, 8.73024e-010, 8.79274e-010,
+ 8.85524e-010, 8.91774e-010, 8.98024e-010, 9.04274e-010, 9.10524e-010, 9.16774e-010,
+ 9.23024e-010, 9.29274e-010, 9.35524e-010, 9.41774e-010, 9.48024e-010, 9.54274e-010,
+ 9.60524e-010, 9.66774e-010, 9.73024e-010, 9.79274e-010, 9.85524e-010, 9.91774e-010,
+ 9.98024e-010, 1.00427e-009, 1.01052e-009, 1.01677e-009, 1.02302e-009, 1.02927e-009,
+ 1.03552e-009, 1.04177e-009, 1.04802e-009, 1.05427e-009, 1.06052e-009, 1.06677e-009,
+ 1.07302e-009, 1.07927e-009, 1.08552e-009, 1.09177e-009, 1.09802e-009, 1.10427e-009,
+ 1.11052e-009, 1.11677e-009, 1.12302e-009, 1.12927e-009, 1.13552e-009, 1.14177e-009,
+ 1.14802e-009, 1.15427e-009, 1.16052e-009, 1.16677e-009, 1.17302e-009, 1.17927e-009,
+ 1.18552e-009, 1.19177e-009, 1.19802e-009, 1.20427e-009, 1.21052e-009, 1.21677e-009,
+ 1.22302e-009, 1.22927e-009, 1.23552e-009, 1.24177e-009, 1.24802e-009, 1.25427e-009,
+ 1.26052e-009, 1.26677e-009, 1.27302e-009, 1.27927e-009, 1.28552e-009, 1.29177e-009,
+ 1.29802e-009, 1.30427e-009, 1.31052e-009, 1.31677e-009, 1.32302e-009, 1.32927e-009,
+ 1.33552e-009, 1.34177e-009, 1.34802e-009, 1.35427e-009, 1.36052e-009, 1.36677e-009,
+ 1.37302e-009, 1.37927e-009, 1.38552e-009, 1.39177e-009, 1.39802e-009, 1.40427e-009,
+ 1.41052e-009, 1.41677e-009, 1.42302e-009, 1.42927e-009, 1.43552e-009, 1.44177e-009,
+ 1.44802e-009, 1.45427e-009, 1.46052e-009, 1.46677e-009)"
+          kdata_1to0_min="(1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 0.994646, 0.993826, 0.993007, 0.992189, 0.980394,
+ 0.978163, 0.975939, 0.973721, 0.97151, 0.945079, 0.939915,
+ 0.93477, 0.929645, 0.924539, 0.91305, 0.907394, 0.901718,
+ 0.896024, 0.890313, 0.817187, 0.80378, 0.790449, 0.777194,
+ 0.764017, 0.726053, 0.710242, 0.694453, 0.67869, 0.55545,
+ 0.528887, 0.502923, 0.477672, 0.452928, 0.441447, 0.417835,
+ 0.394483, 0.371407, 0.348571, 0.281799, 0.255858, 0.230407,
+ 0.20539, 0.180756, 0.195081, 0.173155, 0.151292, 0.129533,
+ 0.107868, 0.118215, 0.0991421, 0.0800503, 0.0609434, 0.0418339,
+ 0.0555166, 0.0392241, 0.0228697, 0.00641968, 0.0495123, 0.0386718,
+ 0.027634, 0.0164357, 0.00508082, 0.0142965, 0.00525532, 0,
+ 0, 0, 0.011854, 0.00700832, 0.00205821, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 5.24679e-005, 0.00025246,
+ 0.000453967, 0.000657004, 0.000861589, 0.00106774, 0.00127547, 0.0014848,
+ 0.00169204, 0.0019002, 0.00210928, 0.00231928, 0.00100161, 0.00100357,
+ 0.00100553, 0.0010075, 0.00100947, 0.00100465, 0.00100577, 0.00100691,
+ 0.00100804, 0.00100918, 0.00101032, 0.00101146, 0.0010126, 0.00101375,
+ 0.00101491, 0.00101366, 0.00101452, 0.00101539, 0.00101627, 0.00101714,
+ 0.00101553, 0.00101612, 0.0010167, 0.00101728, 0.00101787, 0.00101845,
+ 0.00101904, 0.00101962, 0.00102021, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0)"
+          vdata_min="(-0.9, -0.84, -0.78, -0.72, -0.66, -0.6,
+ -0.54, -0.48, -0.42, -0.36, -0.3, -0.24,
+ -0.18, -0.12, -0.06, 0, 0.06, 0.12,
+ 0.18, 0.24, 0.3, 0.36, 0.42, 0.48,
+ 0.54, 0.6, 0.66, 0.72, 0.78, 0.84,
+ 0.9, 0.96, 1.02, 1.08, 1.14, 1.2,
+ 1.26, 1.32, 1.38, 1.44, 1.5, 1.56,
+ 1.62, 1.68, 1.74, 1.8, 1.86, 1.92,
+ 1.98, 2.04, 2.1, 2.16, 2.22, 2.28,
+ 2.34, 2.4, 2.46, 2.52, 2.58, 2.64,
+ 2.7, 2.76, 2.82, 2.88, 2.94, 3,
+ 3.06, 3.12, 3.18, 3.24, 3.3, 3.36,
+ 3.42, 3.48, 3.54, 3.6)"
+          idata_min="(-0.02224, -0.02215, -0.021557, -0.020807, -0.019932, -0.01894,
+ -0.017762, -0.0163597, -0.0146538, -0.0127109, -0.0106332, -0.0085203,
+ -0.0063937, -0.004263, -0.002132, 0, 0.002124, 0.004233,
+ 0.006324, 0.008397, 0.01045, 0.01249, 0.0145, 0.01649,
+ 0.01846, 0.0204, 0.02231, 0.0242, 0.02606, 0.0279,
+ 0.0297, 0.03146, 0.0332, 0.03489, 0.03655, 0.03817,
+ 0.03974, 0.04128, 0.04276, 0.04419, 0.04556, 0.04688,
+ 0.04813, 0.04932, 0.05042, 0.05145, 0.05239, 0.05324,
+ 0.0539998, 0.0546683, 0.0552489, 0.0557519, 0.056186, 0.05657,
+ 0.056897, 0.0572, 0.057457, 0.057706, 0.05793, 0.058132,
+ 0.05833, 0.05856, 0.05869, 0.0588, 0.0591, 0.0592,
+ 0.0593, 0.0594, 0.0596, 0.0598, 0.0599, 0.06,
+ 0.0602, 0.0603, 0.0604, 0.0606)"
+          tdata_0to1_max="(4.96516e-012, 1.23871e-011, 1.9809e-011, 2.7231e-011, 3.46529e-011, 4.20748e-011,
+ 4.94968e-011, 5.69187e-011, 6.43406e-011, 7.17626e-011, 7.91845e-011, 8.66065e-011,
+ 9.40284e-011, 1.0145e-010, 1.08872e-010, 1.16294e-010, 1.23716e-010, 1.31138e-010,
+ 1.3856e-010, 1.45982e-010, 1.53404e-010, 1.60826e-010, 1.68248e-010, 1.7567e-010,
+ 1.83092e-010, 1.90514e-010, 1.97935e-010, 2.05357e-010, 2.12779e-010, 2.20201e-010,
+ 2.27623e-010, 2.35045e-010, 2.42467e-010, 2.49889e-010, 2.57311e-010, 2.64733e-010,
+ 2.72155e-010, 2.79577e-010, 2.86999e-010, 2.94421e-010, 3.01843e-010, 3.09265e-010,
+ 3.16686e-010, 3.24108e-010, 3.3153e-010, 3.38952e-010, 3.46374e-010, 3.53796e-010,
+ 3.61218e-010, 3.6864e-010, 3.76062e-010, 3.83484e-010, 3.90906e-010, 3.98328e-010,
+ 4.0575e-010, 4.13172e-010, 4.20594e-010, 4.28015e-010, 4.35437e-010, 4.42859e-010,
+ 4.50281e-010, 4.57703e-010, 4.65125e-010, 4.72547e-010, 4.79969e-010, 4.87391e-010,
+ 4.94813e-010, 5.02235e-010, 5.09657e-010, 5.17079e-010, 5.24501e-010, 5.31923e-010,
+ 5.39345e-010, 5.46766e-010, 5.54188e-010, 5.6161e-010, 5.69032e-010, 5.76454e-010,
+ 5.83876e-010, 5.91298e-010, 5.9872e-010, 6.06142e-010, 6.13564e-010, 6.20986e-010,
+ 6.28408e-010, 6.3583e-010, 6.43252e-010, 6.50674e-010, 6.58095e-010, 6.65517e-010,
+ 6.72939e-010, 6.80361e-010, 6.87783e-010, 6.95205e-010, 7.02627e-010, 7.10049e-010,
+ 7.17471e-010, 7.24893e-010, 7.32315e-010, 7.39737e-010, 7.47159e-010, 7.54581e-010,
+ 7.62003e-010, 7.69425e-010, 7.76846e-010, 7.84268e-010, 7.9169e-010, 7.99112e-010,
+ 8.06534e-010, 8.13956e-010, 8.21378e-010, 8.288e-010, 8.36222e-010, 8.43644e-010,
+ 8.51066e-010, 8.58488e-010, 8.6591e-010, 8.73332e-010, 8.80754e-010, 8.88175e-010,
+ 8.95597e-010, 9.03019e-010, 9.10441e-010, 9.17863e-010, 9.25285e-010, 9.32707e-010,
+ 9.40129e-010, 9.47551e-010, 9.54973e-010, 9.62395e-010, 9.69817e-010, 9.77239e-010,
+ 9.84661e-010, 9.92083e-010, 9.99505e-010, 1.00693e-009, 1.01435e-009, 1.02177e-009,
+ 1.02919e-009, 1.03661e-009, 1.04404e-009, 1.05146e-009, 1.05888e-009, 1.0663e-009,
+ 1.07372e-009, 1.08115e-009, 1.08857e-009, 1.09599e-009, 1.10341e-009, 1.11083e-009,
+ 1.11826e-009, 1.12568e-009, 1.1331e-009, 1.14052e-009, 1.14794e-009, 1.15537e-009,
+ 1.16279e-009, 1.17021e-009, 1.17763e-009, 1.18505e-009, 1.19247e-009, 1.1999e-009,
+ 1.20732e-009, 1.21474e-009, 1.22216e-009, 1.22958e-009, 1.23701e-009, 1.24443e-009,
+ 1.25185e-009, 1.25927e-009, 1.26669e-009, 1.27412e-009, 1.28154e-009, 1.28896e-009,
+ 1.29638e-009, 1.3038e-009, 1.31123e-009, 1.31865e-009, 1.32607e-009, 1.33349e-009,
+ 1.34091e-009, 1.34834e-009, 1.35576e-009, 1.36318e-009, 1.3706e-009, 1.37802e-009,
+ 1.38545e-009, 1.39287e-009, 1.40029e-009, 1.40771e-009, 1.41513e-009, 1.42255e-009,
+ 1.42998e-009, 1.4374e-009, 1.44482e-009, 1.45224e-009, 1.45966e-009, 1.46709e-009,
+ 1.47451e-009, 1.48193e-009, 1.48935e-009, 1.49677e-009, 1.5042e-009)"
+          kdata_0to1_max="(0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0.00569651, 0.00797394, 0.0101697, 0.0122872, 0.0456626,
+ 0.0510044, 0.0561412, 0.0610819, 0.0899824, 0.0974826, 0.104784,
+ 0.111894, 0.118823, 0.177096, 0.188923, 0.200394, 0.211537,
+ 0.222298, 0.255786, 0.267891, 0.279519, 0.290826, 0.345133,
+ 0.360612, 0.375734, 0.390569, 0.424544, 0.441794, 0.458924,
+ 0.475911, 0.515607, 0.53587, 0.556206, 0.576611, 0.596363,
+ 0.618281, 0.640704, 0.663382, 0.663809, 0.684793, 0.706227,
+ 0.728215, 0.739928, 0.762191, 0.784981, 0.808267, 0.781378,
+ 0.798831, 0.816575, 0.834617, 0.837009, 0.853991, 0.871298,
+ 0.888938, 0.853994, 0.864319, 0.87483, 0.885447, 0.896391,
+ 0.907642, 0.919051, 0.930624, 0.915004, 0.922767, 0.930609,
+ 0.93853, 0.935223, 0.941614, 0.948057, 0.954555, 0.943771,
+ 0.947669, 0.951587, 0.955524, 0.954325, 0.957495, 0.960677,
+ 0.963872, 0.959697, 0.961761, 0.96383, 0.965904, 0.965428,
+ 0.96711, 0.968795, 0.970484, 0.969038, 0.970237, 0.971437,
+ 0.97264, 0.973112, 0.974201, 0.975292, 0.976383, 0.975782,
+ 0.976605, 0.977428, 0.978253, 0.980456, 0.981505, 0.982555,
+ 0.983607, 0.982997, 0.98378, 0.984564, 0.985349, 0.984822,
+ 0.985393, 0.985964, 0.986536, 0.986131, 0.986543, 0.986954,
+ 0.987366, 0.987778, 0.987452, 0.987759, 0.988067, 0.988374,
+ 0.988708, 0.989019, 0.989331, 0.989643, 0.989984, 0.990301,
+ 0.990617, 0.990934, 0.990885, 0.991149, 0.991413, 0.991677,
+ 0.991961, 0.992228, 0.992495, 0.992763, 0.992662, 0.992875,
+ 0.993089, 0.993302, 0.994259, 0.994583, 0.994907, 0.995231,
+ 0.994741, 0.994944, 0.995147, 0.99535, 0.995553, 0.995502,
+ 0.995665, 0.995828, 0.995991, 0.995808, 0.995915, 0.996023,
+ 0.996131, 0.996242, 0.99635, 0.996458, 0.996566, 0.996678,
+ 0.996787, 0.996896, 0.997005, 0.997116, 0.997225, 0.997334,
+ 0.997444, 0.997555, 0.997665, 0.997775, 0.997885, 0.997657,
+ 0.997711, 0.997765, 0.997819, 0.997872, 1)"
+          tdata_1to0_max="(2.10524e-010, 2.16774e-010, 2.23024e-010, 2.29274e-010, 2.35524e-010, 2.41774e-010,
+ 2.48024e-010, 2.54274e-010, 2.60524e-010, 2.66774e-010, 2.73024e-010, 2.79274e-010,
+ 2.85524e-010, 2.91774e-010, 2.98024e-010, 3.04274e-010, 3.10524e-010, 3.16774e-010,
+ 3.23024e-010, 3.29274e-010, 3.35524e-010, 3.41774e-010, 3.48024e-010, 3.54274e-010,
+ 3.60524e-010, 3.66774e-010, 3.73024e-010, 3.79274e-010, 3.85524e-010, 3.91774e-010,
+ 3.98024e-010, 4.04274e-010, 4.10524e-010, 4.16774e-010, 4.23024e-010, 4.29274e-010,
+ 4.35524e-010, 4.41774e-010, 4.48024e-010, 4.54274e-010, 4.60524e-010, 4.66774e-010,
+ 4.73024e-010, 4.79274e-010, 4.85524e-010, 4.91774e-010, 4.98024e-010, 5.04274e-010,
+ 5.10524e-010, 5.16774e-010, 5.23024e-010, 5.29274e-010, 5.35524e-010, 5.41774e-010,
+ 5.48024e-010, 5.54274e-010, 5.60524e-010, 5.66774e-010, 5.73024e-010, 5.79274e-010,
+ 5.85524e-010, 5.91774e-010, 5.98024e-010, 6.04274e-010, 6.10524e-010, 6.16774e-010,
+ 6.23024e-010, 6.29274e-010, 6.35524e-010, 6.41774e-010, 6.48024e-010, 6.54274e-010,
+ 6.60524e-010, 6.66774e-010, 6.73024e-010, 6.79274e-010, 6.85524e-010, 6.91774e-010,
+ 6.98024e-010, 7.04274e-010, 7.10524e-010, 7.16774e-010, 7.23024e-010, 7.29274e-010,
+ 7.35524e-010, 7.41774e-010, 7.48024e-010, 7.54274e-010, 7.60524e-010, 7.66774e-010,
+ 7.73024e-010, 7.79274e-010, 7.85524e-010, 7.91774e-010, 7.98024e-010, 8.04274e-010,
+ 8.10524e-010, 8.16774e-010, 8.23024e-010, 8.29274e-010, 8.35524e-010, 8.41774e-010,
+ 8.48024e-010, 8.54274e-010, 8.60524e-010, 8.66774e-010, 8.73024e-010, 8.79274e-010,
+ 8.85524e-010, 8.91774e-010, 8.98024e-010, 9.04274e-010, 9.10524e-010, 9.16774e-010,
+ 9.23024e-010, 9.29274e-010, 9.35524e-010, 9.41774e-010, 9.48024e-010, 9.54274e-010,
+ 9.60524e-010, 9.66774e-010, 9.73024e-010, 9.79274e-010, 9.85524e-010, 9.91774e-010,
+ 9.98024e-010, 1.00427e-009, 1.01052e-009, 1.01677e-009, 1.02302e-009, 1.02927e-009,
+ 1.03552e-009, 1.04177e-009, 1.04802e-009, 1.05427e-009, 1.06052e-009, 1.06677e-009,
+ 1.07302e-009, 1.07927e-009, 1.08552e-009, 1.09177e-009, 1.09802e-009, 1.10427e-009,
+ 1.11052e-009, 1.11677e-009, 1.12302e-009, 1.12927e-009, 1.13552e-009, 1.14177e-009,
+ 1.14802e-009, 1.15427e-009, 1.16052e-009, 1.16677e-009, 1.17302e-009, 1.17927e-009,
+ 1.18552e-009, 1.19177e-009, 1.19802e-009, 1.20427e-009, 1.21052e-009, 1.21677e-009,
+ 1.22302e-009, 1.22927e-009, 1.23552e-009, 1.24177e-009, 1.24802e-009, 1.25427e-009,
+ 1.26052e-009, 1.26677e-009, 1.27302e-009, 1.27927e-009, 1.28552e-009, 1.29177e-009,
+ 1.29802e-009, 1.30427e-009, 1.31052e-009, 1.31677e-009, 1.32302e-009, 1.32927e-009,
+ 1.33552e-009, 1.34177e-009, 1.34802e-009, 1.35427e-009, 1.36052e-009, 1.36677e-009,
+ 1.37302e-009, 1.37927e-009, 1.38552e-009, 1.39177e-009, 1.39802e-009, 1.40427e-009,
+ 1.41052e-009, 1.41677e-009, 1.42302e-009, 1.42927e-009, 1.43552e-009, 1.44177e-009,
+ 1.44802e-009, 1.45427e-009, 1.46052e-009, 1.46677e-009)"
+          kdata_1to0_max="(1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 0.994646, 0.993826, 0.993007, 0.992189, 0.980394,
+ 0.978163, 0.975939, 0.973721, 0.97151, 0.945079, 0.939915,
+ 0.93477, 0.929645, 0.924539, 0.91305, 0.907394, 0.901718,
+ 0.896024, 0.890313, 0.817187, 0.80378, 0.790449, 0.777194,
+ 0.764017, 0.726053, 0.710242, 0.694453, 0.67869, 0.55545,
+ 0.528887, 0.502923, 0.477672, 0.452928, 0.441447, 0.417835,
+ 0.394483, 0.371407, 0.348571, 0.281799, 0.255858, 0.230407,
+ 0.20539, 0.180756, 0.195081, 0.173155, 0.151292, 0.129533,
+ 0.107868, 0.118215, 0.0991421, 0.0800503, 0.0609434, 0.0418339,
+ 0.0555166, 0.0392241, 0.0228697, 0.00641968, 0.0495123, 0.0386718,
+ 0.027634, 0.0164357, 0.00508082, 0.0142965, 0.00525532, 0,
+ 0, 0, 0.011854, 0.00700832, 0.00205821, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 5.24679e-005, 0.00025246,
+ 0.000453967, 0.000657004, 0.000861589, 0.00106774, 0.00127547, 0.0014848,
+ 0.00169204, 0.0019002, 0.00210928, 0.00231928, 0.00100161, 0.00100357,
+ 0.00100553, 0.0010075, 0.00100947, 0.00100465, 0.00100577, 0.00100691,
+ 0.00100804, 0.00100918, 0.00101032, 0.00101146, 0.0010126, 0.00101375,
+ 0.00101491, 0.00101366, 0.00101452, 0.00101539, 0.00101627, 0.00101714,
+ 0.00101553, 0.00101612, 0.0010167, 0.00101728, 0.00101787, 0.00101845,
+ 0.00101904, 0.00101962, 0.00102021, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0)"
+          vdata_max="(-0.9, -0.84, -0.78, -0.72, -0.66, -0.6,
+ -0.54, -0.48, -0.42, -0.36, -0.3, -0.24,
+ -0.18, -0.12, -0.06, 0, 0.06, 0.12,
+ 0.18, 0.24, 0.3, 0.36, 0.42, 0.48,
+ 0.54, 0.6, 0.66, 0.72, 0.78, 0.84,
+ 0.9, 0.96, 1.02, 1.08, 1.14, 1.2,
+ 1.26, 1.32, 1.38, 1.44, 1.5, 1.56,
+ 1.62, 1.68, 1.74, 1.8, 1.86, 1.92,
+ 1.98, 2.04, 2.1, 2.16, 2.22, 2.28,
+ 2.34, 2.4, 2.46, 2.52, 2.58, 2.64,
+ 2.7, 2.76, 2.82, 2.88, 2.94, 3,
+ 3.06, 3.12, 3.18, 3.24, 3.3, 3.36,
+ 3.42, 3.48, 3.54, 3.6)"
+          idata_max="(-0.02224, -0.02215, -0.021557, -0.020807, -0.019932, -0.01894,
+ -0.017762, -0.0163597, -0.0146538, -0.0127109, -0.0106332, -0.0085203,
+ -0.0063937, -0.004263, -0.002132, 0, 0.002124, 0.004233,
+ 0.006324, 0.008397, 0.01045, 0.01249, 0.0145, 0.01649,
+ 0.01846, 0.0204, 0.02231, 0.0242, 0.02606, 0.0279,
+ 0.0297, 0.03146, 0.0332, 0.03489, 0.03655, 0.03817,
+ 0.03974, 0.04128, 0.04276, 0.04419, 0.04556, 0.04688,
+ 0.04813, 0.04932, 0.05042, 0.05145, 0.05239, 0.05324,
+ 0.0539998, 0.0546683, 0.0552489, 0.0557519, 0.056186, 0.05657,
+ 0.056897, 0.0572, 0.057457, 0.057706, 0.05793, 0.058132,
+ 0.05833, 0.05856, 0.05869, 0.0588, 0.0591, 0.0592,
+ 0.0593, 0.0594, 0.0596, 0.0598, 0.0599, 0.06,
+ 0.0602, 0.0603, 0.0604, 0.0606)"
+ PORT: a_PdRef
+       a_signal
+       d_pulldown_control


*IBIS Pullup tables
Y_PullUp ibis_ktiv(icx_behavioral)
+ GENERIC: corner="ibis_typ"
+          tdata_0to1_typ="(2.10524e-010, 2.16774e-010, 2.23024e-010, 2.29274e-010, 2.35524e-010, 2.41774e-010,
+ 2.48024e-010, 2.54274e-010, 2.60524e-010, 2.66774e-010, 2.73024e-010, 2.79274e-010,
+ 2.85524e-010, 2.91774e-010, 2.98024e-010, 3.04274e-010, 3.10524e-010, 3.16774e-010,
+ 3.23024e-010, 3.29274e-010, 3.35524e-010, 3.41774e-010, 3.48024e-010, 3.54274e-010,
+ 3.60524e-010, 3.66774e-010, 3.73024e-010, 3.79274e-010, 3.85524e-010, 3.91774e-010,
+ 3.98024e-010, 4.04274e-010, 4.10524e-010, 4.16774e-010, 4.23024e-010, 4.29274e-010,
+ 4.35524e-010, 4.41774e-010, 4.48024e-010, 4.54274e-010, 4.60524e-010, 4.66774e-010,
+ 4.73024e-010, 4.79274e-010, 4.85524e-010, 4.91774e-010, 4.98024e-010, 5.04274e-010,
+ 5.10524e-010, 5.16774e-010, 5.23024e-010, 5.29274e-010, 5.35524e-010, 5.41774e-010,
+ 5.48024e-010, 5.54274e-010, 5.60524e-010, 5.66774e-010, 5.73024e-010, 5.79274e-010,
+ 5.85524e-010, 5.91774e-010, 5.98024e-010, 6.04274e-010, 6.10524e-010, 6.16774e-010,
+ 6.23024e-010, 6.29274e-010, 6.35524e-010, 6.41774e-010, 6.48024e-010, 6.54274e-010,
+ 6.60524e-010, 6.66774e-010, 6.73024e-010, 6.79274e-010, 6.85524e-010, 6.91774e-010,
+ 6.98024e-010, 7.04274e-010, 7.10524e-010, 7.16774e-010, 7.23024e-010, 7.29274e-010,
+ 7.35524e-010, 7.41774e-010, 7.48024e-010, 7.54274e-010, 7.60524e-010, 7.66774e-010,
+ 7.73024e-010, 7.79274e-010, 7.85524e-010, 7.91774e-010, 7.98024e-010, 8.04274e-010,
+ 8.10524e-010, 8.16774e-010, 8.23024e-010, 8.29274e-010, 8.35524e-010, 8.41774e-010,
+ 8.48024e-010, 8.54274e-010, 8.60524e-010, 8.66774e-010, 8.73024e-010, 8.79274e-010,
+ 8.85524e-010, 8.91774e-010, 8.98024e-010, 9.04274e-010, 9.10524e-010, 9.16774e-010,
+ 9.23024e-010, 9.29274e-010, 9.35524e-010, 9.41774e-010, 9.48024e-010, 9.54274e-010,
+ 9.60524e-010, 9.66774e-010, 9.73024e-010, 9.79274e-010, 9.85524e-010, 9.91774e-010,
+ 9.98024e-010, 1.00427e-009, 1.01052e-009, 1.01677e-009, 1.02302e-009, 1.02927e-009,
+ 1.03552e-009, 1.04177e-009, 1.04802e-009, 1.05427e-009, 1.06052e-009, 1.06677e-009,
+ 1.07302e-009, 1.07927e-009, 1.08552e-009, 1.09177e-009, 1.09802e-009, 1.10427e-009,
+ 1.11052e-009, 1.11677e-009, 1.12302e-009, 1.12927e-009, 1.13552e-009, 1.14177e-009,
+ 1.14802e-009, 1.15427e-009, 1.16052e-009, 1.16677e-009, 1.17302e-009, 1.17927e-009,
+ 1.18552e-009, 1.19177e-009, 1.19802e-009, 1.20427e-009, 1.21052e-009, 1.21677e-009,
+ 1.22302e-009, 1.22927e-009, 1.23552e-009, 1.24177e-009, 1.24802e-009, 1.25427e-009,
+ 1.26052e-009, 1.26677e-009, 1.27302e-009, 1.27927e-009, 1.28552e-009, 1.29177e-009,
+ 1.29802e-009, 1.30427e-009, 1.31052e-009, 1.31677e-009, 1.32302e-009, 1.32927e-009,
+ 1.33552e-009, 1.34177e-009, 1.34802e-009, 1.35427e-009, 1.36052e-009, 1.36677e-009,
+ 1.37302e-009, 1.37927e-009, 1.38552e-009, 1.39177e-009, 1.39802e-009, 1.40427e-009,
+ 1.41052e-009, 1.41677e-009, 1.42302e-009, 1.42927e-009, 1.43552e-009, 1.44177e-009,
+ 1.44802e-009, 1.45427e-009, 1.46052e-009, 1.46677e-009)"
+          kdata_0to1_typ="(0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0.00146725, 0.00341046,
+ 0.00534272, 0.00726409, 0.00917463, 0.0413965, 0.0474324, 0.0534458,
+ 0.0594367, 0.065405, 0.085689, 0.0931554, 0.100517, 0.107774,
+ 0.114927, 0.16011, 0.171528, 0.18277, 0.193835, 0.200159,
+ 0.20938, 0.218257, 0.226811, 0.235034, 0.290475, 0.303465,
+ 0.316046, 0.328223, 0.340061, 0.345863, 0.355782, 0.365274,
+ 0.374341, 0.382936, 0.438353, 0.451142, 0.463458, 0.475401,
+ 0.486927, 0.509469, 0.521916, 0.533981, 0.545671, 0.557063,
+ 0.567685, 0.578964, 0.590052, 0.600794, 0.644498, 0.659791,
+ 0.675007, 0.690258, 0.705564, 0.674914, 0.685555, 0.69628,
+ 0.706936, 0.717519, 0.761797, 0.777244, 0.792863, 0.808664,
+ 0.824648, 0.780955, 0.790848, 0.800805, 0.810826, 0.820911,
+ 0.848496, 0.861157, 0.87413, 0.887286, 0.850574, 0.857796,
+ 0.865072, 0.8724, 0.879781, 0.896427, 0.905214, 0.914119,
+ 0.923188, 0.932356, 0.910489, 0.916065, 0.921681, 0.927338,
+ 0.933037, 0.938777, 0.944559, 0.950384, 0.956253, 0.962165,
+ 0.94564, 0.94896, 0.952293, 0.955641, 0.956699, 0.959752,
+ 0.962816, 0.965892, 0.968979, 0.961439, 0.963203, 0.964971,
+ 0.966742, 0.968517, 0.970296, 0.972079, 0.973866, 0.975663,
+ 0.977469, 0.975513, 0.97687, 0.978229, 0.97959, 0.980954,
+ 0.978447, 0.979357, 0.980267, 0.981179, 0.982091, 0.983005,
+ 0.983919, 0.984835, 0.985751, 0.984188, 0.984769, 0.985349,
+ 0.98593, 0.986511, 0.985933, 0.986392, 0.986852, 0.987312,
+ 0.987772, 0.988232, 0.988693, 0.989154, 0.989615, 0.990076,
+ 0.992494, 0.993188, 0.993882, 0.994578, 0.993943, 0.994464,
+ 0.994986, 0.995509, 0.996031, 0.996554, 0.997078, 0.993287,
+ 0.993287, 0.993287, 0.993287, 0.993287, 0.993287, 0.993287,
+ 0.993287, 0.993287, 0.996843, 0.997308, 0.997774, 0.99824,
+ 0.998706, 0.995519, 0.995519, 0.995519, 0.995519, 0.995519,
+ 0.995519, 0.995519, 0.995519, 0.995519, 0.995519, 0.999359,
+ 0.999826, 1, 1, 1)"
+          tdata_1to0_typ="(4.96516e-012, 1.23871e-011, 1.9809e-011, 2.7231e-011, 3.46529e-011, 4.20748e-011,
+ 4.94968e-011, 5.69187e-011, 6.43406e-011, 7.17626e-011, 7.91845e-011, 8.66065e-011,
+ 9.40284e-011, 1.0145e-010, 1.08872e-010, 1.16294e-010, 1.23716e-010, 1.31138e-010,
+ 1.3856e-010, 1.45982e-010, 1.53404e-010, 1.60826e-010, 1.68248e-010, 1.7567e-010,
+ 1.83092e-010, 1.90514e-010, 1.97935e-010, 2.05357e-010, 2.12779e-010, 2.20201e-010,
+ 2.27623e-010, 2.35045e-010, 2.42467e-010, 2.49889e-010, 2.57311e-010, 2.64733e-010,
+ 2.72155e-010, 2.79577e-010, 2.86999e-010, 2.94421e-010, 3.01843e-010, 3.09265e-010,
+ 3.16686e-010, 3.24108e-010, 3.3153e-010, 3.38952e-010, 3.46374e-010, 3.53796e-010,
+ 3.61218e-010, 3.6864e-010, 3.76062e-010, 3.83484e-010, 3.90906e-010, 3.98328e-010,
+ 4.0575e-010, 4.13172e-010, 4.20594e-010, 4.28015e-010, 4.35437e-010, 4.42859e-010,
+ 4.50281e-010, 4.57703e-010, 4.65125e-010, 4.72547e-010, 4.79969e-010, 4.87391e-010,
+ 4.94813e-010, 5.02235e-010, 5.09657e-010, 5.17079e-010, 5.24501e-010, 5.31923e-010,
+ 5.39345e-010, 5.46766e-010, 5.54188e-010, 5.6161e-010, 5.69032e-010, 5.76454e-010,
+ 5.83876e-010, 5.91298e-010, 5.9872e-010, 6.06142e-010, 6.13564e-010, 6.20986e-010,
+ 6.28408e-010, 6.3583e-010, 6.43252e-010, 6.50674e-010, 6.58095e-010, 6.65517e-010,
+ 6.72939e-010, 6.80361e-010, 6.87783e-010, 6.95205e-010, 7.02627e-010, 7.10049e-010,
+ 7.17471e-010, 7.24893e-010, 7.32315e-010, 7.39737e-010, 7.47159e-010, 7.54581e-010,
+ 7.62003e-010, 7.69425e-010, 7.76846e-010, 7.84268e-010, 7.9169e-010, 7.99112e-010,
+ 8.06534e-010, 8.13956e-010, 8.21378e-010, 8.288e-010, 8.36222e-010, 8.43644e-010,
+ 8.51066e-010, 8.58488e-010, 8.6591e-010, 8.73332e-010, 8.80754e-010, 8.88175e-010,
+ 8.95597e-010, 9.03019e-010, 9.10441e-010, 9.17863e-010, 9.25285e-010, 9.32707e-010,
+ 9.40129e-010, 9.47551e-010, 9.54973e-010, 9.62395e-010, 9.69817e-010, 9.77239e-010,
+ 9.84661e-010, 9.92083e-010, 9.99505e-010, 1.00693e-009, 1.01435e-009, 1.02177e-009,
+ 1.02919e-009, 1.03661e-009, 1.04404e-009, 1.05146e-009, 1.05888e-009, 1.0663e-009,
+ 1.07372e-009, 1.08115e-009, 1.08857e-009, 1.09599e-009, 1.10341e-009, 1.11083e-009,
+ 1.11826e-009, 1.12568e-009, 1.1331e-009, 1.14052e-009, 1.14794e-009, 1.15537e-009,
+ 1.16279e-009, 1.17021e-009, 1.17763e-009, 1.18505e-009, 1.19247e-009, 1.1999e-009,
+ 1.20732e-009, 1.21474e-009, 1.22216e-009, 1.22958e-009, 1.23701e-009, 1.24443e-009,
+ 1.25185e-009, 1.25927e-009, 1.26669e-009, 1.27412e-009, 1.28154e-009, 1.28896e-009,
+ 1.29638e-009, 1.3038e-009, 1.31123e-009, 1.31865e-009, 1.32607e-009, 1.33349e-009,
+ 1.34091e-009, 1.34834e-009, 1.35576e-009, 1.36318e-009, 1.3706e-009, 1.37802e-009,
+ 1.38545e-009, 1.39287e-009, 1.40029e-009, 1.40771e-009, 1.41513e-009, 1.42255e-009,
+ 1.42998e-009, 1.4374e-009, 1.44482e-009, 1.45224e-009, 1.45966e-009, 1.46709e-009,
+ 1.47451e-009, 1.48193e-009, 1.48935e-009, 1.49677e-009, 1.5042e-009)"
+          kdata_1to0_typ="(1, 0.9946, 0.993782, 0.992965, 0.992149, 0.980948,
+ 0.978649, 0.976358, 0.974075, 0.956583, 0.952217, 0.947877,
+ 0.943565, 0.920627, 0.913868, 0.907172, 0.900537, 0.850466,
+ 0.838511, 0.826752, 0.815184, 0.749376, 0.731983, 0.715011,
+ 0.698446, 0.604929, 0.581536, 0.55887, 0.536954, 0.477789,
+ 0.45349, 0.429952, 0.407104, 0.434402, 0.416594, 0.398965,
+ 0.381542, 0.36439, 0.303333, 0.281306, 0.25942, 0.237733,
+ 0.21619, 0.183612, 0.160801, 0.138016, 0.115368, 0.136067,
+ 0.116059, 0.0958237, 0.075428, 0.100249, 0.0833551, 0.0661689,
+ 0.0486857, 0.066046, 0.0512897, 0.0361615, 0.0206773, 0.0532476,
+ 0.0427263, 0.0319095, 0.0207627, 0.0285438, 0.0193926, 0.00999358,
+ 0.000344576, 0.0236224, 0.0180178, 0.0122248, 0.00623936, 0.0090203,
+ 0.00420322, 0, 0, 0.00573283, 0.00297215, 0.000148583,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0.00114683, 0.00129392, 0.00144257,
+ 0.00159282, 0.00141581, 0.00151547, 0.00161599, 0.00171737, 0.00146279,
+ 0.00150711, 0.00155165, 0.00159642, 0.00140687, 0.00141363, 0.00142041,
+ 0.00142722, 0.00134165, 0.0013333, 0.00132493, 0.00131654, 0.00120915,
+ 0.00118425, 0.0011593, 0.00113429, 0.00108017, 0.00105026, 0.0010203,
+ 0.00099029, 0.000928789, 0.000893374, 0.000857909, 0.000822395, 0.000795697,
+ 0.00076166, 0.000727587, 0.000693478, 0.000671278, 0.000639119, 0.000606918,
+ 0.000574673, 0.00056284, 0.000534127, 0.000505386, 0.000476616, 0.000471733,
+ 0.000447148, 0.000422546, 0.000397926, 0.000392937, 0.000371789, 0.00035063,
+ 0.000329459, 0.000308278, 0.000313783, 0.000296645, 0.000279499, 0.000262348,
+ 0.000262702, 0.000248213, 0.000233718, 0.000219218, 0.000224494, 0.000213027,
+ 0.000201555, 0.000190079, 0.000189821, 0.000180079, 0.000170333, 0.000160584,
+ 0.00016385, 0.000156126, 0.0001484, 0.000140672, 0.000139903, 0.000133266,
+ 0.000126627, 0.000119986, 0.000106635, 9.89244e-005, 9.12101e-005, 8.34927e-005,
+ 9.49625e-005, 9.03043e-005, 8.5645e-005, 8.09844e-005, 7.63226e-005, 7.89374e-005,
+ 7.55122e-005, 7.20863e-005, 6.86597e-005, 6.83e-005, 6.53987e-005, 6.2497e-005,
+ 5.95949e-005, 5.85277e-005, 5.59417e-005, 5.33553e-005, 5.07685e-005, 5.03451e-005,
+ 4.8134e-005, 4.59225e-005, 4.37108e-005, 4.28391e-005, 4.08617e-005, 3.8884e-005,
+ 3.69061e-005, 3.65148e-005, 3.48166e-005, 3.31181e-005, 3.14194e-005, 3.07619e-005,
+ 2.92486e-005, 2.77352e-005, 2.62217e-005, 2.47081e-005, 0)"
+          vdata_typ="(-1.8, -1.32, -1.26, -1.2, -1.14, -1.08,
+ -1.02, -0.96, -0.9, -0.84, -0.78, -0.72,
+ -0.66, -0.6, -0.54, -0.48, -0.42, -0.36,
+ -0.3, -0.24, -0.18, -0.12, -0.06, 0,
+ 0.06, 0.12, 0.18, 0.24, 0.3, 0.36,
+ 0.42, 0.48, 0.54, 0.6, 0.66, 0.72,
+ 0.78, 0.84, 0.9, 0.96, 1.02, 1.08,
+ 1.14, 1.2, 1.26, 1.32, 1.38, 1.44,
+ 1.5, 1.56, 1.62, 1.68, 1.74, 1.8,
+ 1.86, 1.92, 1.98, 2.04, 2.1, 2.16,
+ 2.22, 2.28, 2.34, 2.4, 2.46, 2.52,
+ 2.58)"
+          idata_typ="(-0.0263, -0.0263, -0.0262, -0.0259, -0.0255, -0.0249,
+ -0.02429, -0.0236, -0.02286, -0.022052, -0.0212, -0.020266,
+ -0.019257, -0.01814, -0.016897, -0.01546, -0.013806, -0.0119419,
+ -0.0099739, -0.0079753, -0.0059738, -0.003976, -0.001985, 2.09e-010,
+ 0.001974, 0.003933, 0.005876, 0.007803, 0.009712, 0.0116,
+ 0.01348, 0.01533, 0.01716, 0.01897, 0.02075, 0.02251,
+ 0.02425, 0.02596, 0.02764, 0.02929, 0.03091, 0.0325,
+ 0.03406, 0.03558, 0.03706, 0.03851, 0.03991, 0.04127,
+ 0.04258, 0.04385, 0.04506, 0.04622, 0.04732, 0.04836,
+ 0.04933, 0.05024, 0.0510797, 0.0518673, 0.0525732, 0.0532309,
+ 0.0538338, 0.0543897, 0.054902, 0.05539, 0.055832, 0.056247,
+ 0.056527)"
+          tdata_0to1_min="(2.10524e-010, 2.16774e-010, 2.23024e-010, 2.29274e-010, 2.35524e-010, 2.41774e-010,
+ 2.48024e-010, 2.54274e-010, 2.60524e-010, 2.66774e-010, 2.73024e-010, 2.79274e-010,
+ 2.85524e-010, 2.91774e-010, 2.98024e-010, 3.04274e-010, 3.10524e-010, 3.16774e-010,
+ 3.23024e-010, 3.29274e-010, 3.35524e-010, 3.41774e-010, 3.48024e-010, 3.54274e-010,
+ 3.60524e-010, 3.66774e-010, 3.73024e-010, 3.79274e-010, 3.85524e-010, 3.91774e-010,
+ 3.98024e-010, 4.04274e-010, 4.10524e-010, 4.16774e-010, 4.23024e-010, 4.29274e-010,
+ 4.35524e-010, 4.41774e-010, 4.48024e-010, 4.54274e-010, 4.60524e-010, 4.66774e-010,
+ 4.73024e-010, 4.79274e-010, 4.85524e-010, 4.91774e-010, 4.98024e-010, 5.04274e-010,
+ 5.10524e-010, 5.16774e-010, 5.23024e-010, 5.29274e-010, 5.35524e-010, 5.41774e-010,
+ 5.48024e-010, 5.54274e-010, 5.60524e-010, 5.66774e-010, 5.73024e-010, 5.79274e-010,
+ 5.85524e-010, 5.91774e-010, 5.98024e-010, 6.04274e-010, 6.10524e-010, 6.16774e-010,
+ 6.23024e-010, 6.29274e-010, 6.35524e-010, 6.41774e-010, 6.48024e-010, 6.54274e-010,
+ 6.60524e-010, 6.66774e-010, 6.73024e-010, 6.79274e-010, 6.85524e-010, 6.91774e-010,
+ 6.98024e-010, 7.04274e-010, 7.10524e-010, 7.16774e-010, 7.23024e-010, 7.29274e-010,
+ 7.35524e-010, 7.41774e-010, 7.48024e-010, 7.54274e-010, 7.60524e-010, 7.66774e-010,
+ 7.73024e-010, 7.79274e-010, 7.85524e-010, 7.91774e-010, 7.98024e-010, 8.04274e-010,
+ 8.10524e-010, 8.16774e-010, 8.23024e-010, 8.29274e-010, 8.35524e-010, 8.41774e-010,
+ 8.48024e-010, 8.54274e-010, 8.60524e-010, 8.66774e-010, 8.73024e-010, 8.79274e-010,
+ 8.85524e-010, 8.91774e-010, 8.98024e-010, 9.04274e-010, 9.10524e-010, 9.16774e-010,
+ 9.23024e-010, 9.29274e-010, 9.35524e-010, 9.41774e-010, 9.48024e-010, 9.54274e-010,
+ 9.60524e-010, 9.66774e-010, 9.73024e-010, 9.79274e-010, 9.85524e-010, 9.91774e-010,
+ 9.98024e-010, 1.00427e-009, 1.01052e-009, 1.01677e-009, 1.02302e-009, 1.02927e-009,
+ 1.03552e-009, 1.04177e-009, 1.04802e-009, 1.05427e-009, 1.06052e-009, 1.06677e-009,
+ 1.07302e-009, 1.07927e-009, 1.08552e-009, 1.09177e-009, 1.09802e-009, 1.10427e-009,
+ 1.11052e-009, 1.11677e-009, 1.12302e-009, 1.12927e-009, 1.13552e-009, 1.14177e-009,
+ 1.14802e-009, 1.15427e-009, 1.16052e-009, 1.16677e-009, 1.17302e-009, 1.17927e-009,
+ 1.18552e-009, 1.19177e-009, 1.19802e-009, 1.20427e-009, 1.21052e-009, 1.21677e-009,
+ 1.22302e-009, 1.22927e-009, 1.23552e-009, 1.24177e-009, 1.24802e-009, 1.25427e-009,
+ 1.26052e-009, 1.26677e-009, 1.27302e-009, 1.27927e-009, 1.28552e-009, 1.29177e-009,
+ 1.29802e-009, 1.30427e-009, 1.31052e-009, 1.31677e-009, 1.32302e-009, 1.32927e-009,
+ 1.33552e-009, 1.34177e-009, 1.34802e-009, 1.35427e-009, 1.36052e-009, 1.36677e-009,
+ 1.37302e-009, 1.37927e-009, 1.38552e-009, 1.39177e-009, 1.39802e-009, 1.40427e-009,
+ 1.41052e-009, 1.41677e-009, 1.42302e-009, 1.42927e-009, 1.43552e-009, 1.44177e-009,
+ 1.44802e-009, 1.45427e-009, 1.46052e-009, 1.46677e-009)"
+          kdata_0to1_min="(0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0.00146725, 0.00341046,
+ 0.00534272, 0.00726409, 0.00917463, 0.0413965, 0.0474324, 0.0534458,
+ 0.0594367, 0.065405, 0.085689, 0.0931554, 0.100517, 0.107774,
+ 0.114927, 0.16011, 0.171528, 0.18277, 0.193835, 0.200159,
+ 0.20938, 0.218257, 0.226811, 0.235034, 0.290475, 0.303465,
+ 0.316046, 0.328223, 0.340061, 0.345863, 0.355782, 0.365274,
+ 0.374341, 0.382936, 0.438353, 0.451142, 0.463458, 0.475401,
+ 0.486927, 0.509469, 0.521916, 0.533981, 0.545671, 0.557063,
+ 0.567685, 0.578964, 0.590052, 0.600794, 0.644498, 0.659791,
+ 0.675007, 0.690258, 0.705564, 0.674914, 0.685555, 0.69628,
+ 0.706936, 0.717519, 0.761797, 0.777244, 0.792863, 0.808664,
+ 0.824648, 0.780955, 0.790848, 0.800805, 0.810826, 0.820911,
+ 0.848496, 0.861157, 0.87413, 0.887286, 0.850574, 0.857796,
+ 0.865072, 0.8724, 0.879781, 0.896427, 0.905214, 0.914119,
+ 0.923188, 0.932356, 0.910489, 0.916065, 0.921681, 0.927338,
+ 0.933037, 0.938777, 0.944559, 0.950384, 0.956253, 0.962165,
+ 0.94564, 0.94896, 0.952293, 0.955641, 0.956699, 0.959752,
+ 0.962816, 0.965892, 0.968979, 0.961439, 0.963203, 0.964971,
+ 0.966742, 0.968517, 0.970296, 0.972079, 0.973866, 0.975663,
+ 0.977469, 0.975513, 0.97687, 0.978229, 0.97959, 0.980954,
+ 0.978447, 0.979357, 0.980267, 0.981179, 0.982091, 0.983005,
+ 0.983919, 0.984835, 0.985751, 0.984188, 0.984769, 0.985349,
+ 0.98593, 0.986511, 0.985933, 0.986392, 0.986852, 0.987312,
+ 0.987772, 0.988232, 0.988693, 0.989154, 0.989615, 0.990076,
+ 0.992494, 0.993188, 0.993882, 0.994578, 0.993943, 0.994464,
+ 0.994986, 0.995509, 0.996031, 0.996554, 0.997078, 0.993287,
+ 0.993287, 0.993287, 0.993287, 0.993287, 0.993287, 0.993287,
+ 0.993287, 0.993287, 0.996843, 0.997308, 0.997774, 0.99824,
+ 0.998706, 0.995519, 0.995519, 0.995519, 0.995519, 0.995519,
+ 0.995519, 0.995519, 0.995519, 0.995519, 0.995519, 0.999359,
+ 0.999826, 1, 1, 1)"
+          tdata_1to0_min="(4.96516e-012, 1.23871e-011, 1.9809e-011, 2.7231e-011, 3.46529e-011, 4.20748e-011,
+ 4.94968e-011, 5.69187e-011, 6.43406e-011, 7.17626e-011, 7.91845e-011, 8.66065e-011,
+ 9.40284e-011, 1.0145e-010, 1.08872e-010, 1.16294e-010, 1.23716e-010, 1.31138e-010,
+ 1.3856e-010, 1.45982e-010, 1.53404e-010, 1.60826e-010, 1.68248e-010, 1.7567e-010,
+ 1.83092e-010, 1.90514e-010, 1.97935e-010, 2.05357e-010, 2.12779e-010, 2.20201e-010,
+ 2.27623e-010, 2.35045e-010, 2.42467e-010, 2.49889e-010, 2.57311e-010, 2.64733e-010,
+ 2.72155e-010, 2.79577e-010, 2.86999e-010, 2.94421e-010, 3.01843e-010, 3.09265e-010,
+ 3.16686e-010, 3.24108e-010, 3.3153e-010, 3.38952e-010, 3.46374e-010, 3.53796e-010,
+ 3.61218e-010, 3.6864e-010, 3.76062e-010, 3.83484e-010, 3.90906e-010, 3.98328e-010,
+ 4.0575e-010, 4.13172e-010, 4.20594e-010, 4.28015e-010, 4.35437e-010, 4.42859e-010,
+ 4.50281e-010, 4.57703e-010, 4.65125e-010, 4.72547e-010, 4.79969e-010, 4.87391e-010,
+ 4.94813e-010, 5.02235e-010, 5.09657e-010, 5.17079e-010, 5.24501e-010, 5.31923e-010,
+ 5.39345e-010, 5.46766e-010, 5.54188e-010, 5.6161e-010, 5.69032e-010, 5.76454e-010,
+ 5.83876e-010, 5.91298e-010, 5.9872e-010, 6.06142e-010, 6.13564e-010, 6.20986e-010,
+ 6.28408e-010, 6.3583e-010, 6.43252e-010, 6.50674e-010, 6.58095e-010, 6.65517e-010,
+ 6.72939e-010, 6.80361e-010, 6.87783e-010, 6.95205e-010, 7.02627e-010, 7.10049e-010,
+ 7.17471e-010, 7.24893e-010, 7.32315e-010, 7.39737e-010, 7.47159e-010, 7.54581e-010,
+ 7.62003e-010, 7.69425e-010, 7.76846e-010, 7.84268e-010, 7.9169e-010, 7.99112e-010,
+ 8.06534e-010, 8.13956e-010, 8.21378e-010, 8.288e-010, 8.36222e-010, 8.43644e-010,
+ 8.51066e-010, 8.58488e-010, 8.6591e-010, 8.73332e-010, 8.80754e-010, 8.88175e-010,
+ 8.95597e-010, 9.03019e-010, 9.10441e-010, 9.17863e-010, 9.25285e-010, 9.32707e-010,
+ 9.40129e-010, 9.47551e-010, 9.54973e-010, 9.62395e-010, 9.69817e-010, 9.77239e-010,
+ 9.84661e-010, 9.92083e-010, 9.99505e-010, 1.00693e-009, 1.01435e-009, 1.02177e-009,
+ 1.02919e-009, 1.03661e-009, 1.04404e-009, 1.05146e-009, 1.05888e-009, 1.0663e-009,
+ 1.07372e-009, 1.08115e-009, 1.08857e-009, 1.09599e-009, 1.10341e-009, 1.11083e-009,
+ 1.11826e-009, 1.12568e-009, 1.1331e-009, 1.14052e-009, 1.14794e-009, 1.15537e-009,
+ 1.16279e-009, 1.17021e-009, 1.17763e-009, 1.18505e-009, 1.19247e-009, 1.1999e-009,
+ 1.20732e-009, 1.21474e-009, 1.22216e-009, 1.22958e-009, 1.23701e-009, 1.24443e-009,
+ 1.25185e-009, 1.25927e-009, 1.26669e-009, 1.27412e-009, 1.28154e-009, 1.28896e-009,
+ 1.29638e-009, 1.3038e-009, 1.31123e-009, 1.31865e-009, 1.32607e-009, 1.33349e-009,
+ 1.34091e-009, 1.34834e-009, 1.35576e-009, 1.36318e-009, 1.3706e-009, 1.37802e-009,
+ 1.38545e-009, 1.39287e-009, 1.40029e-009, 1.40771e-009, 1.41513e-009, 1.42255e-009,
+ 1.42998e-009, 1.4374e-009, 1.44482e-009, 1.45224e-009, 1.45966e-009, 1.46709e-009,
+ 1.47451e-009, 1.48193e-009, 1.48935e-009, 1.49677e-009, 1.5042e-009)"
+          kdata_1to0_min="(1, 0.9946, 0.993782, 0.992965, 0.992149, 0.980948,
+ 0.978649, 0.976358, 0.974075, 0.956583, 0.952217, 0.947877,
+ 0.943565, 0.920627, 0.913868, 0.907172, 0.900537, 0.850466,
+ 0.838511, 0.826752, 0.815184, 0.749376, 0.731983, 0.715011,
+ 0.698446, 0.604929, 0.581536, 0.55887, 0.536954, 0.477789,
+ 0.45349, 0.429952, 0.407104, 0.434402, 0.416594, 0.398965,
+ 0.381542, 0.36439, 0.303333, 0.281306, 0.25942, 0.237733,
+ 0.21619, 0.183612, 0.160801, 0.138016, 0.115368, 0.136067,
+ 0.116059, 0.0958237, 0.075428, 0.100249, 0.0833551, 0.0661689,
+ 0.0486857, 0.066046, 0.0512897, 0.0361615, 0.0206773, 0.0532476,
+ 0.0427263, 0.0319095, 0.0207627, 0.0285438, 0.0193926, 0.00999358,
+ 0.000344576, 0.0236224, 0.0180178, 0.0122248, 0.00623936, 0.0090203,
+ 0.00420322, 0, 0, 0.00573283, 0.00297215, 0.000148583,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0.00114683, 0.00129392, 0.00144257,
+ 0.00159282, 0.00141581, 0.00151547, 0.00161599, 0.00171737, 0.00146279,
+ 0.00150711, 0.00155165, 0.00159642, 0.00140687, 0.00141363, 0.00142041,
+ 0.00142722, 0.00134165, 0.0013333, 0.00132493, 0.00131654, 0.00120915,
+ 0.00118425, 0.0011593, 0.00113429, 0.00108017, 0.00105026, 0.0010203,
+ 0.00099029, 0.000928789, 0.000893374, 0.000857909, 0.000822395, 0.000795697,
+ 0.00076166, 0.000727587, 0.000693478, 0.000671278, 0.000639119, 0.000606918,
+ 0.000574673, 0.00056284, 0.000534127, 0.000505386, 0.000476616, 0.000471733,
+ 0.000447148, 0.000422546, 0.000397926, 0.000392937, 0.000371789, 0.00035063,
+ 0.000329459, 0.000308278, 0.000313783, 0.000296645, 0.000279499, 0.000262348,
+ 0.000262702, 0.000248213, 0.000233718, 0.000219218, 0.000224494, 0.000213027,
+ 0.000201555, 0.000190079, 0.000189821, 0.000180079, 0.000170333, 0.000160584,
+ 0.00016385, 0.000156126, 0.0001484, 0.000140672, 0.000139903, 0.000133266,
+ 0.000126627, 0.000119986, 0.000106635, 9.89244e-005, 9.12101e-005, 8.34927e-005,
+ 9.49625e-005, 9.03043e-005, 8.5645e-005, 8.09844e-005, 7.63226e-005, 7.89374e-005,
+ 7.55122e-005, 7.20863e-005, 6.86597e-005, 6.83e-005, 6.53987e-005, 6.2497e-005,
+ 5.95949e-005, 5.85277e-005, 5.59417e-005, 5.33553e-005, 5.07685e-005, 5.03451e-005,
+ 4.8134e-005, 4.59225e-005, 4.37108e-005, 4.28391e-005, 4.08617e-005, 3.8884e-005,
+ 3.69061e-005, 3.65148e-005, 3.48166e-005, 3.31181e-005, 3.14194e-005, 3.07619e-005,
+ 2.92486e-005, 2.77352e-005, 2.62217e-005, 2.47081e-005, 0)"
+          vdata_min="(-1.8, -1.32, -1.26, -1.2, -1.14, -1.08,
+ -1.02, -0.96, -0.9, -0.84, -0.78, -0.72,
+ -0.66, -0.6, -0.54, -0.48, -0.42, -0.36,
+ -0.3, -0.24, -0.18, -0.12, -0.06, 0,
+ 0.06, 0.12, 0.18, 0.24, 0.3, 0.36,
+ 0.42, 0.48, 0.54, 0.6, 0.66, 0.72,
+ 0.78, 0.84, 0.9, 0.96, 1.02, 1.08,
+ 1.14, 1.2, 1.26, 1.32, 1.38, 1.44,
+ 1.5, 1.56, 1.62, 1.68, 1.74, 1.8,
+ 1.86, 1.92, 1.98, 2.04, 2.1, 2.16,
+ 2.22, 2.28, 2.34, 2.4, 2.46, 2.52,
+ 2.58)"
+          idata_min="(-0.0263, -0.0263, -0.0262, -0.0259, -0.0255, -0.0249,
+ -0.02429, -0.0236, -0.02286, -0.022052, -0.0212, -0.020266,
+ -0.019257, -0.01814, -0.016897, -0.01546, -0.013806, -0.0119419,
+ -0.0099739, -0.0079753, -0.0059738, -0.003976, -0.001985, 2.09e-010,
+ 0.001974, 0.003933, 0.005876, 0.007803, 0.009712, 0.0116,
+ 0.01348, 0.01533, 0.01716, 0.01897, 0.02075, 0.02251,
+ 0.02425, 0.02596, 0.02764, 0.02929, 0.03091, 0.0325,
+ 0.03406, 0.03558, 0.03706, 0.03851, 0.03991, 0.04127,
+ 0.04258, 0.04385, 0.04506, 0.04622, 0.04732, 0.04836,
+ 0.04933, 0.05024, 0.0510797, 0.0518673, 0.0525732, 0.0532309,
+ 0.0538338, 0.0543897, 0.054902, 0.05539, 0.055832, 0.056247,
+ 0.056527)"
+          tdata_0to1_max="(2.10524e-010, 2.16774e-010, 2.23024e-010, 2.29274e-010, 2.35524e-010, 2.41774e-010,
+ 2.48024e-010, 2.54274e-010, 2.60524e-010, 2.66774e-010, 2.73024e-010, 2.79274e-010,
+ 2.85524e-010, 2.91774e-010, 2.98024e-010, 3.04274e-010, 3.10524e-010, 3.16774e-010,
+ 3.23024e-010, 3.29274e-010, 3.35524e-010, 3.41774e-010, 3.48024e-010, 3.54274e-010,
+ 3.60524e-010, 3.66774e-010, 3.73024e-010, 3.79274e-010, 3.85524e-010, 3.91774e-010,
+ 3.98024e-010, 4.04274e-010, 4.10524e-010, 4.16774e-010, 4.23024e-010, 4.29274e-010,
+ 4.35524e-010, 4.41774e-010, 4.48024e-010, 4.54274e-010, 4.60524e-010, 4.66774e-010,
+ 4.73024e-010, 4.79274e-010, 4.85524e-010, 4.91774e-010, 4.98024e-010, 5.04274e-010,
+ 5.10524e-010, 5.16774e-010, 5.23024e-010, 5.29274e-010, 5.35524e-010, 5.41774e-010,
+ 5.48024e-010, 5.54274e-010, 5.60524e-010, 5.66774e-010, 5.73024e-010, 5.79274e-010,
+ 5.85524e-010, 5.91774e-010, 5.98024e-010, 6.04274e-010, 6.10524e-010, 6.16774e-010,
+ 6.23024e-010, 6.29274e-010, 6.35524e-010, 6.41774e-010, 6.48024e-010, 6.54274e-010,
+ 6.60524e-010, 6.66774e-010, 6.73024e-010, 6.79274e-010, 6.85524e-010, 6.91774e-010,
+ 6.98024e-010, 7.04274e-010, 7.10524e-010, 7.16774e-010, 7.23024e-010, 7.29274e-010,
+ 7.35524e-010, 7.41774e-010, 7.48024e-010, 7.54274e-010, 7.60524e-010, 7.66774e-010,
+ 7.73024e-010, 7.79274e-010, 7.85524e-010, 7.91774e-010, 7.98024e-010, 8.04274e-010,
+ 8.10524e-010, 8.16774e-010, 8.23024e-010, 8.29274e-010, 8.35524e-010, 8.41774e-010,
+ 8.48024e-010, 8.54274e-010, 8.60524e-010, 8.66774e-010, 8.73024e-010, 8.79274e-010,
+ 8.85524e-010, 8.91774e-010, 8.98024e-010, 9.04274e-010, 9.10524e-010, 9.16774e-010,
+ 9.23024e-010, 9.29274e-010, 9.35524e-010, 9.41774e-010, 9.48024e-010, 9.54274e-010,
+ 9.60524e-010, 9.66774e-010, 9.73024e-010, 9.79274e-010, 9.85524e-010, 9.91774e-010,
+ 9.98024e-010, 1.00427e-009, 1.01052e-009, 1.01677e-009, 1.02302e-009, 1.02927e-009,
+ 1.03552e-009, 1.04177e-009, 1.04802e-009, 1.05427e-009, 1.06052e-009, 1.06677e-009,
+ 1.07302e-009, 1.07927e-009, 1.08552e-009, 1.09177e-009, 1.09802e-009, 1.10427e-009,
+ 1.11052e-009, 1.11677e-009, 1.12302e-009, 1.12927e-009, 1.13552e-009, 1.14177e-009,
+ 1.14802e-009, 1.15427e-009, 1.16052e-009, 1.16677e-009, 1.17302e-009, 1.17927e-009,
+ 1.18552e-009, 1.19177e-009, 1.19802e-009, 1.20427e-009, 1.21052e-009, 1.21677e-009,
+ 1.22302e-009, 1.22927e-009, 1.23552e-009, 1.24177e-009, 1.24802e-009, 1.25427e-009,
+ 1.26052e-009, 1.26677e-009, 1.27302e-009, 1.27927e-009, 1.28552e-009, 1.29177e-009,
+ 1.29802e-009, 1.30427e-009, 1.31052e-009, 1.31677e-009, 1.32302e-009, 1.32927e-009,
+ 1.33552e-009, 1.34177e-009, 1.34802e-009, 1.35427e-009, 1.36052e-009, 1.36677e-009,
+ 1.37302e-009, 1.37927e-009, 1.38552e-009, 1.39177e-009, 1.39802e-009, 1.40427e-009,
+ 1.41052e-009, 1.41677e-009, 1.42302e-009, 1.42927e-009, 1.43552e-009, 1.44177e-009,
+ 1.44802e-009, 1.45427e-009, 1.46052e-009, 1.46677e-009)"
+          kdata_0to1_max="(0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0.00146725, 0.00341046,
+ 0.00534272, 0.00726409, 0.00917463, 0.0413965, 0.0474324, 0.0534458,
+ 0.0594367, 0.065405, 0.085689, 0.0931554, 0.100517, 0.107774,
+ 0.114927, 0.16011, 0.171528, 0.18277, 0.193835, 0.200159,
+ 0.20938, 0.218257, 0.226811, 0.235034, 0.290475, 0.303465,
+ 0.316046, 0.328223, 0.340061, 0.345863, 0.355782, 0.365274,
+ 0.374341, 0.382936, 0.438353, 0.451142, 0.463458, 0.475401,
+ 0.486927, 0.509469, 0.521916, 0.533981, 0.545671, 0.557063,
+ 0.567685, 0.578964, 0.590052, 0.600794, 0.644498, 0.659791,
+ 0.675007, 0.690258, 0.705564, 0.674914, 0.685555, 0.69628,
+ 0.706936, 0.717519, 0.761797, 0.777244, 0.792863, 0.808664,
+ 0.824648, 0.780955, 0.790848, 0.800805, 0.810826, 0.820911,
+ 0.848496, 0.861157, 0.87413, 0.887286, 0.850574, 0.857796,
+ 0.865072, 0.8724, 0.879781, 0.896427, 0.905214, 0.914119,
+ 0.923188, 0.932356, 0.910489, 0.916065, 0.921681, 0.927338,
+ 0.933037, 0.938777, 0.944559, 0.950384, 0.956253, 0.962165,
+ 0.94564, 0.94896, 0.952293, 0.955641, 0.956699, 0.959752,
+ 0.962816, 0.965892, 0.968979, 0.961439, 0.963203, 0.964971,
+ 0.966742, 0.968517, 0.970296, 0.972079, 0.973866, 0.975663,
+ 0.977469, 0.975513, 0.97687, 0.978229, 0.97959, 0.980954,
+ 0.978447, 0.979357, 0.980267, 0.981179, 0.982091, 0.983005,
+ 0.983919, 0.984835, 0.985751, 0.984188, 0.984769, 0.985349,
+ 0.98593, 0.986511, 0.985933, 0.986392, 0.986852, 0.987312,
+ 0.987772, 0.988232, 0.988693, 0.989154, 0.989615, 0.990076,
+ 0.992494, 0.993188, 0.993882, 0.994578, 0.993943, 0.994464,
+ 0.994986, 0.995509, 0.996031, 0.996554, 0.997078, 0.993287,
+ 0.993287, 0.993287, 0.993287, 0.993287, 0.993287, 0.993287,
+ 0.993287, 0.993287, 0.996843, 0.997308, 0.997774, 0.99824,
+ 0.998706, 0.995519, 0.995519, 0.995519, 0.995519, 0.995519,
+ 0.995519, 0.995519, 0.995519, 0.995519, 0.995519, 0.999359,
+ 0.999826, 1, 1, 1)"
+          tdata_1to0_max="(4.96516e-012, 1.23871e-011, 1.9809e-011, 2.7231e-011, 3.46529e-011, 4.20748e-011,
+ 4.94968e-011, 5.69187e-011, 6.43406e-011, 7.17626e-011, 7.91845e-011, 8.66065e-011,
+ 9.40284e-011, 1.0145e-010, 1.08872e-010, 1.16294e-010, 1.23716e-010, 1.31138e-010,
+ 1.3856e-010, 1.45982e-010, 1.53404e-010, 1.60826e-010, 1.68248e-010, 1.7567e-010,
+ 1.83092e-010, 1.90514e-010, 1.97935e-010, 2.05357e-010, 2.12779e-010, 2.20201e-010,
+ 2.27623e-010, 2.35045e-010, 2.42467e-010, 2.49889e-010, 2.57311e-010, 2.64733e-010,
+ 2.72155e-010, 2.79577e-010, 2.86999e-010, 2.94421e-010, 3.01843e-010, 3.09265e-010,
+ 3.16686e-010, 3.24108e-010, 3.3153e-010, 3.38952e-010, 3.46374e-010, 3.53796e-010,
+ 3.61218e-010, 3.6864e-010, 3.76062e-010, 3.83484e-010, 3.90906e-010, 3.98328e-010,
+ 4.0575e-010, 4.13172e-010, 4.20594e-010, 4.28015e-010, 4.35437e-010, 4.42859e-010,
+ 4.50281e-010, 4.57703e-010, 4.65125e-010, 4.72547e-010, 4.79969e-010, 4.87391e-010,
+ 4.94813e-010, 5.02235e-010, 5.09657e-010, 5.17079e-010, 5.24501e-010, 5.31923e-010,
+ 5.39345e-010, 5.46766e-010, 5.54188e-010, 5.6161e-010, 5.69032e-010, 5.76454e-010,
+ 5.83876e-010, 5.91298e-010, 5.9872e-010, 6.06142e-010, 6.13564e-010, 6.20986e-010,
+ 6.28408e-010, 6.3583e-010, 6.43252e-010, 6.50674e-010, 6.58095e-010, 6.65517e-010,
+ 6.72939e-010, 6.80361e-010, 6.87783e-010, 6.95205e-010, 7.02627e-010, 7.10049e-010,
+ 7.17471e-010, 7.24893e-010, 7.32315e-010, 7.39737e-010, 7.47159e-010, 7.54581e-010,
+ 7.62003e-010, 7.69425e-010, 7.76846e-010, 7.84268e-010, 7.9169e-010, 7.99112e-010,
+ 8.06534e-010, 8.13956e-010, 8.21378e-010, 8.288e-010, 8.36222e-010, 8.43644e-010,
+ 8.51066e-010, 8.58488e-010, 8.6591e-010, 8.73332e-010, 8.80754e-010, 8.88175e-010,
+ 8.95597e-010, 9.03019e-010, 9.10441e-010, 9.17863e-010, 9.25285e-010, 9.32707e-010,
+ 9.40129e-010, 9.47551e-010, 9.54973e-010, 9.62395e-010, 9.69817e-010, 9.77239e-010,
+ 9.84661e-010, 9.92083e-010, 9.99505e-010, 1.00693e-009, 1.01435e-009, 1.02177e-009,
+ 1.02919e-009, 1.03661e-009, 1.04404e-009, 1.05146e-009, 1.05888e-009, 1.0663e-009,
+ 1.07372e-009, 1.08115e-009, 1.08857e-009, 1.09599e-009, 1.10341e-009, 1.11083e-009,
+ 1.11826e-009, 1.12568e-009, 1.1331e-009, 1.14052e-009, 1.14794e-009, 1.15537e-009,
+ 1.16279e-009, 1.17021e-009, 1.17763e-009, 1.18505e-009, 1.19247e-009, 1.1999e-009,
+ 1.20732e-009, 1.21474e-009, 1.22216e-009, 1.22958e-009, 1.23701e-009, 1.24443e-009,
+ 1.25185e-009, 1.25927e-009, 1.26669e-009, 1.27412e-009, 1.28154e-009, 1.28896e-009,
+ 1.29638e-009, 1.3038e-009, 1.31123e-009, 1.31865e-009, 1.32607e-009, 1.33349e-009,
+ 1.34091e-009, 1.34834e-009, 1.35576e-009, 1.36318e-009, 1.3706e-009, 1.37802e-009,
+ 1.38545e-009, 1.39287e-009, 1.40029e-009, 1.40771e-009, 1.41513e-009, 1.42255e-009,
+ 1.42998e-009, 1.4374e-009, 1.44482e-009, 1.45224e-009, 1.45966e-009, 1.46709e-009,
+ 1.47451e-009, 1.48193e-009, 1.48935e-009, 1.49677e-009, 1.5042e-009)"
+          kdata_1to0_max="(1, 0.9946, 0.993782, 0.992965, 0.992149, 0.980948,
+ 0.978649, 0.976358, 0.974075, 0.956583, 0.952217, 0.947877,
+ 0.943565, 0.920627, 0.913868, 0.907172, 0.900537, 0.850466,
+ 0.838511, 0.826752, 0.815184, 0.749376, 0.731983, 0.715011,
+ 0.698446, 0.604929, 0.581536, 0.55887, 0.536954, 0.477789,
+ 0.45349, 0.429952, 0.407104, 0.434402, 0.416594, 0.398965,
+ 0.381542, 0.36439, 0.303333, 0.281306, 0.25942, 0.237733,
+ 0.21619, 0.183612, 0.160801, 0.138016, 0.115368, 0.136067,
+ 0.116059, 0.0958237, 0.075428, 0.100249, 0.0833551, 0.0661689,
+ 0.0486857, 0.066046, 0.0512897, 0.0361615, 0.0206773, 0.0532476,
+ 0.0427263, 0.0319095, 0.0207627, 0.0285438, 0.0193926, 0.00999358,
+ 0.000344576, 0.0236224, 0.0180178, 0.0122248, 0.00623936, 0.0090203,
+ 0.00420322, 0, 0, 0.00573283, 0.00297215, 0.000148583,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0.00114683, 0.00129392, 0.00144257,
+ 0.00159282, 0.00141581, 0.00151547, 0.00161599, 0.00171737, 0.00146279,
+ 0.00150711, 0.00155165, 0.00159642, 0.00140687, 0.00141363, 0.00142041,
+ 0.00142722, 0.00134165, 0.0013333, 0.00132493, 0.00131654, 0.00120915,
+ 0.00118425, 0.0011593, 0.00113429, 0.00108017, 0.00105026, 0.0010203,
+ 0.00099029, 0.000928789, 0.000893374, 0.000857909, 0.000822395, 0.000795697,
+ 0.00076166, 0.000727587, 0.000693478, 0.000671278, 0.000639119, 0.000606918,
+ 0.000574673, 0.00056284, 0.000534127, 0.000505386, 0.000476616, 0.000471733,
+ 0.000447148, 0.000422546, 0.000397926, 0.000392937, 0.000371789, 0.00035063,
+ 0.000329459, 0.000308278, 0.000313783, 0.000296645, 0.000279499, 0.000262348,
+ 0.000262702, 0.000248213, 0.000233718, 0.000219218, 0.000224494, 0.000213027,
+ 0.000201555, 0.000190079, 0.000189821, 0.000180079, 0.000170333, 0.000160584,
+ 0.00016385, 0.000156126, 0.0001484, 0.000140672, 0.000139903, 0.000133266,
+ 0.000126627, 0.000119986, 0.000106635, 9.89244e-005, 9.12101e-005, 8.34927e-005,
+ 9.49625e-005, 9.03043e-005, 8.5645e-005, 8.09844e-005, 7.63226e-005, 7.89374e-005,
+ 7.55122e-005, 7.20863e-005, 6.86597e-005, 6.83e-005, 6.53987e-005, 6.2497e-005,
+ 5.95949e-005, 5.85277e-005, 5.59417e-005, 5.33553e-005, 5.07685e-005, 5.03451e-005,
+ 4.8134e-005, 4.59225e-005, 4.37108e-005, 4.28391e-005, 4.08617e-005, 3.8884e-005,
+ 3.69061e-005, 3.65148e-005, 3.48166e-005, 3.31181e-005, 3.14194e-005, 3.07619e-005,
+ 2.92486e-005, 2.77352e-005, 2.62217e-005, 2.47081e-005, 0)"
+          vdata_max="(-1.8, -1.32, -1.26, -1.2, -1.14, -1.08,
+ -1.02, -0.96, -0.9, -0.84, -0.78, -0.72,
+ -0.66, -0.6, -0.54, -0.48, -0.42, -0.36,
+ -0.3, -0.24, -0.18, -0.12, -0.06, 0,
+ 0.06, 0.12, 0.18, 0.24, 0.3, 0.36,
+ 0.42, 0.48, 0.54, 0.6, 0.66, 0.72,
+ 0.78, 0.84, 0.9, 0.96, 1.02, 1.08,
+ 1.14, 1.2, 1.26, 1.32, 1.38, 1.44,
+ 1.5, 1.56, 1.62, 1.68, 1.74, 1.8,
+ 1.86, 1.92, 1.98, 2.04, 2.1, 2.16,
+ 2.22, 2.28, 2.34, 2.4, 2.46, 2.52,
+ 2.58)"
+          idata_max="(-0.0263, -0.0263, -0.0262, -0.0259, -0.0255, -0.0249,
+ -0.02429, -0.0236, -0.02286, -0.022052, -0.0212, -0.020266,
+ -0.019257, -0.01814, -0.016897, -0.01546, -0.013806, -0.0119419,
+ -0.0099739, -0.0079753, -0.0059738, -0.003976, -0.001985, 2.09e-010,
+ 0.001974, 0.003933, 0.005876, 0.007803, 0.009712, 0.0116,
+ 0.01348, 0.01533, 0.01716, 0.01897, 0.02075, 0.02251,
+ 0.02425, 0.02596, 0.02764, 0.02929, 0.03091, 0.0325,
+ 0.03406, 0.03558, 0.03706, 0.03851, 0.03991, 0.04127,
+ 0.04258, 0.04385, 0.04506, 0.04622, 0.04732, 0.04836,
+ 0.04933, 0.05024, 0.0510797, 0.0518673, 0.0525732, 0.0532309,
+ 0.0538338, 0.0543897, 0.054902, 0.05539, 0.055832, 0.056247,
+ 0.056527)"
+ PORT: a_signal
+       a_PuRef
+       d_pullup_control

.model ibis_ktiv(icx_behavioral) MACRO LANG=VHDLAMS LIB=icxbase
.ends MODEL_U1_AM10

