***** AD8011 SPICE model       Rev A SMR/ADI 9-30-97

* Copyright 1997 by Analog Devices, Inc.

* Refer to "README.DOC" file for License Statement.  Use of this model
* indicates your acceptance with the terms and provisions in the License Statement.

* This model will give typical performance characteristics
* for the following parameters;

*     closed loop gain and phase vs bandwidth
*     output current and voltage limiting
*     offset voltage (is static, will not vary with vcm)
*     ibias (again, is static, will not vary with vcm)
*     slew rate and step response performance
*     (slew rate is based on 10-90% of step response)
*     current on output will be reflected to the supplies 
*     vnoise, referred to the input
*     inoise, referred to the input

*     distortion is not characterized

* Node assignments
*                non-inverting input
*                | inverting input
*                | | positive supply
*                | | |  negative supply
*                | | |  |  output
*                | | |  |  |
.SUBCKT AD8011an 1 2 99 50 28

* input stage *

q1 50 3 5 qp1
q2 99 5 4 qn1
q3 99 3 6 qn1
q4 50 6 4 qp1
i1 99 5 0.26e-3
i2 6 50 0.26e-3
cin1 1 98 1e-12
cin2 2 98 2.3e-12
v1 4 2 0

* input error sources *

eos 3 1 poly(1) 20 98 2e-3 1
fbn 2 98 poly(1) vnoise3 5e-6 1e-3
fbp 1 98 poly(1) vnoise3 5e-6 1e-3

* gain stage *

f1 98 7 poly(1) v1 0 1 0 100
rgain 7 98 1.3e6
cgain 7 98 1.5e-12
dcl1 7 8 d1
dcl2 9 7 d1
vcl1 99 8 1.54
vcl2 9 50 1.54

gcm 98 7 poly(2) 98 0 30 0 0 1e-5 1e-5

* second pole *

epole 14 98 7 98 1
rpole 14 15 1
cpole 15 98 0.4e-9

* reference stage *

eref 98 0 poly(2) 99 0 50 0 0 0.5 0.5 

ecmref 30 0 poly(2) 1 0 2 0 0 0.5 0.5

* vnoise stage *

rnoise1 19 98 10.6e-3
vnoise1 19 98 0
vnoise2 21 98 0.53
dnoise1 21 19 dn

fnoise1 20 98 vnoise1 1
rnoise2 20 98 1

* inoise stage *

rnoise3 22 98 0.46e-3
vnoise3 22 98 0
vnoise4 24 98 0.6
dnoise2 24 22 dn

fnoise2 23 98 vnoise3 1
rnoise4 23 98 1

* buffer stage *

gbuf 98 13 15 98 1e-2
rbuf 98 13 1e2

* output current reflected to supplies *

fcurr 98 40 voc 1
vcur1 26 98 0
vcur2 98 27 0
dcur1 40 26 d1
dcur2 27 40 d1

* output stage *

vo1 99 90 0
vo2 91 50 0
fout1 0 99 poly(2) vo1 vcur1 -9.27e-3 1 -1
fout2 50 0 poly(2) vo2 vcur2 -9.27e-3 1 -1 
gout1 90 10 13 99 0.1
gout2 91 10 13 50 0.1
rout1 10 90 10
rout2 10 91 10
voc 10 28 0
rout3 28 98 1e6
dcl3 13 11 d1
dcl4 12 13 d1
vcl3 11 10 -0.64
vcl4 10 12 -0.64


.model qp1 pnp(kf=1e-30)
.model qn1 npn(kf=1e-30)
.model d1  d(af=0 kf=1e-30)
.model dn  d(af=1 kf=1e-8)
.ends ad8011an
