* OP421G SPICE Macro-model                 5/91, Rev. A
*                                           JCB / PMI
*
*
* Copyright 1991 by Analog Devices, Inc.
*
* Refer to "README.DOC" file for License Statement.  Use of this model
* indicates your acceptance with the terms and provisions in the License Statement.
*
* Node assignments
*                non-inverting input
*                | inverting input
*                | | positive supply
*                | | |  negative supply
*                | | |  |  output
*                | | |  |  |
.SUBCKT OP421G   1 2 99 50 31
*
* INPUT STAGE & POLE AT 2.8 MEGHZ
*
R1    2  3     5E11
R2    1  3     5E11
R3    5 50     5.16K
R4    6 50     5.16K
CIN   1  2     2E-12
C2    5  6     5.51E-12
I1    99 4     10UA
IOS   1  2     10E-9
EOS   9  1     POLY(1)  24 27  4000E-6  1
Q1    5  2  4  QX
Q2    6  9  4  QX
*
EREF  98 0    27  0  1
*
* FIRST GAIN STAGE
*
R5   10 98     1E6
G1   98 10     5  6  23.1E-6
D1   10 11     DX
D2   12 10     DX
E1   99 11     POLY(1) 99 27 -0.4 1
E2   12 50     POLY(1) 27 50 -0.4 1
*
* GAIN STAGE & DOMINANT POLE AT 9.2 HZ
*
R6   13 98     0.865E9
C3   13 98     20E-12
G2   98 13     10  27   5E-6
V1   99 14     1.7
V2   15 50     1.4
D3   13 14     DX
D4   15 13     DX
*
* POLE AT 3.0 MEGHZ
*
R9   16 98     1E6
C5   16 98     53.1E-15
G3   98 16     13 27  1E-6
*
* POLE AT 3.0 MEGHZ
*
R15  17 98     1E6
C7   17 98     53.1E-15
G10  98 17     16 27  1E-6
**
* COMMON-MODE GAIN NETWORK WITH ZERO AT 30 KHZ
*
R7   24 98     1
R8   23 24     1E6
C4   23 24     5.3E-12
E4   98 23     3  27  100
*
* POLE AT 3.0 MEGHZ
*
R14  25 98     1E6
C6   25 98     53.1E-15
G9   98 25     17 27  1E-6
*
* OUTPUT STAGE
*
ISY  99 50     1040E-6
R10  27 99     33.3E3
R11  27 50     33.3E3
R12  30 99     450
R13  30 50     450
L1   30 31     1E-8
G4   28 50     25 30  2.22E-3
G5   29 50     30 25  2.22E-3
G6   30 99     99 25  2.22E-3
G7   50 30     25 50  2.22E-3
D5   99 28     DX
D6   99 29     DX
D7   50 28     DY
D8   50 29     DY
D9   25 33     DX
V3   33 30     1.7
D10  32 25     DX
V4   30 32     1.7
*
* MODELS USED
*
.MODEL QX PNP(BF=62.5)
.MODEL DX   D(IS=1E-15)
.MODEL DY   D(IS=1E-15 BV=50)
.ENDS
