*AD8002A SPICE Macro Model          11/95, Rev. A
*                                         RFD/ADS
*  
* Copyright 1995 by Analog Devices, Inc.
*
* This version of the AD8002 model simulates the typical 
* parameters of the 'A' grade part.  
*
* This model was developed using the +/-5V specifications.
*
* Refer to the "README.DOC" file for License Statement.  Use of this model
* indicates your acceptance with the terms and provisions in the License  
* Statement.
*
* Node assignments
*               Non-inverting input
*               | Inverting input
*               | | Positive supply
*               | | | Negative supply
*               | | | | Output
*               | | | | |
.SUBCKT AD8002A 3 2 7 4 6 
*
****** INPUT STAGE ******
*
Q1 7 9 10 QN
Q2 4 9 11 QP
Q3 14 11 15 QN
Q4 16 10 15 QP
I1 10 4 DC 2.568e-4 
I2 7 11 DC 2.568e-4 
D1 17 14 DX 
D2 16 18 DX 
V2 18 4 DC -4.41135e-2 
V1 7 17 DC -4.41135e-2 
R1 14 7 1E3 
R2 4 16 1E3 
CS1 7 2 .235e-12 
CS2 2 4 .235e-12 
CIN 3 4 1.5E-12 
LIN- 15 2 .9e-9 
GB1 7 3 POLY(1) 3 100 (3e-6,0.2e-6)
GB2 7 2 POLY(1) 3 100 (5e-6,0.3e-6)
EOS 3 9 POLY(1) 100 23 (2E-3,1)
*
****** GAIN STAGE  ********
*
V3 7 20 DC 2.4 
V4 21 4 DC 2.4 
R3 100 19 9e5 
C1 19 100 6.1e-13 
D3 19 20 DX 
D4 21 19 DX 
G1 100 19 POLY(1) 7 14 (0.0,1E-3)
G2 19 100 POLY(1) 16 4 (0.0,1E-3)
EREF 100 0 POLY(2) (7,0) (4,0) (0,0.5,0.5)
*
****** CMRR STAGE ******
*
CCM 22 23 4.56424e-13 
RCM2 100 23 1 
RCM1 23 22 1e4 
ECM 22 100 POLY(1) 100 3 (0.0,31.668)
*
****** POLE STAGE AT   ******
*
C3 100 24 2.273642e-16 
R5 24 100 1e6 
G4 100 24 POLY(1) 19 100 (0.0,1E-6)
*
****** POLE STAGE AT   ******
*
C4 25 100 3.978877e-17 
R6 25 100 1e6 
G5 100 25 POLY(1) 24 100 (0.0,1E-6)
* 
****** OUTPUT STAGE ****** 
* 
RO1 33 7 21.4 
RO2 4 33 21.4 
VW 25 30 DC 0 
VSC1 31 33 DC .58 
VSC2 33 32 DC .58 
LO 33 6 2e-9 
DSC2 32 30 DX 
DSC1 30 31 DX 
GO1 33 7 POLY(1) 7 30 (0.0,4.6728972e-2)
GO2 4 33 POLY(1) 30 4 (0.0,4.6728972e-2)
*
VSY1 36 100 DC 0 
VSY2 100 37 DC 0 
DSY1 35 36 DX 
DSY2 37 35 DX 
FSY 7 4 POLY(2) VSY1 VSY2 (4.7326E-3,1,1)
GSY 100 35 33 30 4.6728972E-2
*
.MODEL QN NPN(BF=100 IS=1E-15)
.MODEL QP PNP(BF=100 IS=1E-15)
.MODEL DX D(IS=1E-15)
.ENDS AD8002A
