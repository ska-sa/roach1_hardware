*AD8001A SPICE Macro Model       9/94, Rev. A
* AAG/ADSC
*
* Copyright 1994 by Analog Devices, Inc.
*
* Refer to the "README.DOC" file for License Statement.  Use of this model
* indicates your acceptance with the terms and provisions in the License
* Statement
*
* Node assignments
*               Non-inverting input
*               | Inverting input
*               | | Positive supply
*               | | | Negative supply
*               | | | | Output
*               | | | | |
.SUBCKT AD8001A 3 2 7 4 6
*
* INPUT STAGE
*
CIN 3 4 1.5E-12
GB1 7 3 POLY(1) 3 100 (3E-6,0.2E-6)
EOS 9 3 POLY(1) 23 100 (2E-3,1)
Q1 7 9 10 QN
I1 10 4 DC 2.568E-4
I2 7 11 DC 2.568E-4
Q2 4 9 11 QP
R1 7 14 1E3
V1 7 17 DC 6.96561E-2
D1 17 14 DX
Q3 14 11 15 QN
Q4 16 10 15 QP
R2 16 4 1E3
D2 16 18 DX
V2 18 4 DC 6.96561E-2
LIN- 15 2 0.1E-9
GB2 7 2 POLY(1) 3 100 (5E-6,0.3E-6)
CS1 7 2 0.03E-12
CS2 2 4 0.03E-12
*
* GAIN STAGE AND DOMINANT POLE AT 230 kHz
*
EREF 100 0 POLY(2) (7,0) (4,0) (0,0.5,0.5)
G1 100 19 7 14 1E-3
G2 19 100 16 4 1E-3
R3 19 100 1.24E6
C1 19 100 5.580468E-13
V3 7 20 DC 2.3747
D3 19 20 DX
D4 21 19 DX
V4 21 4 DC 2.3747
*
* COMMON-MODE REJECTION NETWORK WITH ZERO AT 22 MHz
*
ECM 100 22 3 100 19.95
RCM1 22 23 1E4
CCM 22 23 7.2343E-13
RCM2 23 100 1
*
* POLE AT 800 MHz
*
G4 100 24 19 100 1E-6
R5 24 100 1E6
C3 24 100 1.9894368E-16
*
* POLE AT 4 GHz
*
G5 100 25 24 100 1E-6
R6 25 100 1E6
C4 25 100 3.9788736E-17
*
* OUTPUT STAGE
*
VW 25 30 DC 0
*
FSY 7 4 POLY(2) VSY1 VSY2 (4.2326E-3,1,1)
GSY 100 35 33 30 4.6728972E-2
DSY1 35 36 DX
VSY1 36 100 DC 0
DSY2 37 35 DX
VSY2 100 37 DC 0
DSC1 30 31 DX
VSC1 31 33 DC 0.62526
DSC2 32 30 DX
VSC2 33 32 DC 0.62526
GO1 33 7 7 30 4.6728972E-2
RO1 7 33 21.4
GO2 4 33 30 4 4.6728972E-2
RO2 33 4 21.4
LO 33 6 7E-9
*
.MODEL QN NPN(BF=100 IS=1E-15)
.MODEL QP PNP(BF=100 IS=1E-15)
.MODEL DX D(IS=1E-15)
*
.ENDS AD8001A
