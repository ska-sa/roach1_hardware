* OP220F SPICE Macro-model                 9/91, Rev. A
*                                           JCB / PMI
*
* This version of the OP-220 model simulates the worst case 
* parameters of the 'F' grade.  The worst case parameters
* used correspond to those in the data sheet.
*
* Copyright 1991 by Analog Devices, Inc.
*
* Refer to "README.DOC" file for License Statement.  Use of this model
* indicates your acceptance with the terms and provisions in the License Statement.
*
* Node assignments
*               non-inverting input
*               | inverting input
*               | | positive supply
*               | | |  negative supply
*               | | |  |  output
*               | | |  |  |
.SUBCKT OP220F  1 2 99 50 30
*
* INPUT STAGE & POLE AT 1.5 MEGHZ
*
R1    2  3     5E11
R2    1  3     5E11
R3    5 50     5.16K
R4    6 50     5.16K
CIN   1  2     4E-12
C2    5  6     15.42E-12
I1    99 4     10UA
IOS   1  2     1.0E-9
EOS   9  1     POLY(1)  24 27  300E-6  1
Q1    5  2  4  QX
Q2    6  9  4  QX
*
EREF  98 0    27  0  1
*
* FIRST GAIN STAGE
*
R5   10 98     1E6
G1   98 10     5  6  50.27E-6
D1   10 11     DX
D2   12 10     DX
E1   99 11     POLY(1) 99 27 -1.475 1
E2   12 50     POLY(1) 27 50 -1.475 1
*
* GAIN STAGE & DOMINANT POLE AT 0.2 HZ
*
R6   13 98     3.98E9
C3   13 98     200E-12
G2   98 13     10 27  5E-6
V1   99 14     1.0
V2   15 50     1.0
D3   13 14     DX
D4   15 13     DX
*
* COMMON-MODE GAIN NETWORK WITH ZERO AT 632 HZ
*
R7   24 98     1
R8   23 24     1E6
C4   23 24     0.252E-9
E4   98 23     3  27  31.6
*
* POLE AT 600 KHZ
*
R9   25 98     1E6
C5   25 98     265E-15
G3   98 25     13 27  1E-6
*
* OUTPUT STAGE
*
ISY  99 50     43.6E-6
R10  27 99     568E3
R11  27 50     568E3
R12  30 99     2000
R13  30 50     2000
G4   28 50     25 30  0.5E-3
G5   29 50     30 25  0.5E-3
G6   30 99     99 25  0.5E-3
G7   50 30     25 50  0.5E-3
D5   99 28     DX
D6   99 29     DX
D7   50 28     DY
D8   50 29     DY
D9   25 31     DX
V3   31 30     3.1
D10  32 25     DX
V4   30 32     0.5
*
* MODELS USED
*
.MODEL QX PNP(BF=200)
.MODEL DX   D(IS=1E-15)
.MODEL DY   D(IS=1E-15 BV=50)
.ENDS
