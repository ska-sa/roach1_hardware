* AD600J SPICE Macro-model              Rev. A, 2/93
*                                       ARG / PMI
*
* This version of the AD600 model simulates the worst case 
* parameters of the 'J' grade.  The worst case parameters
* used correspond to those in the data sheet.
*
* Copyright 1993 by Analog Devices
*
* Refer to "README.DOC" file for License Statement.  Use of
* this model indicates your acceptance of the terms and pro-
* visions in the License Statement.
*
* Node assignments
*                input HI
*                |  input LO
*                |  |  positive supply
*                |  |  |  negative supply
*                |  |  |  |  output
*                |  |  |  |  |  control HI
*                |  |  |  |  |  |  control LO
*                |  |  |  |  |  |  |  gate input
*                |  |  |  |  |  |  |  |  output common
*                |  |  |  |  |  |  |  |  |
.SUBCKT AD600J   3  2  99 50 48 40 41 70 12
*
* INPUT STAGE
*
Q1A  1    3    21   QN
Q1B  4    5    21   QN
Q2A  1    14   22   QN
Q2B  4    5    22   QN
Q3A  1    15   23   QN
Q3B  4    5    23   QN
Q4A  1    16   24   QN
Q4B  4    5    24   QN
Q5A  1    17   25   QN
Q5B  4    5    25   QN
Q6A  1    18   26   QN
Q6B  4    5    26   QN
Q7A  1    19   27   QN
Q7B  4    5    27   QN
Q8A  1    20   28   QN
Q8B  4    5    28   QN
RT   3    2    500
RL1  3    14   62.5
RL2  14   2    125
RL3  14   15   62.5
RL4  15   2    125
RL5  15   16   62.5
RL6  16   2    125
RL7  16   17   62.5
RL8  17   2    125
RL9  17   18   62.5
RL10 18   2    125
RL11 18   19   62.5
RL12 19   2    125
RL13 19   20   62.5
RL14 20   2    62.5
EOS  11   5    POLY(2) (12,2) (38,98) 420E-6 8.84E-3 8.84E-3
RCM  12   98   40E3
IB1  99   7    400E-6
IB2  99   29   200E-6
IB3  99   30   200E-6
IB4  99   31   200E-6
IB5  99   32   200E-6
IB6  99   33   200E-6
IB7  99   34   200E-6
IB8  99   13   400E-6
E1   7    50   POLY(1) (40,41) 2.8 2.4
E2   13   50   POLY(1) (41,40) 2.8 2.4
RB1  7    29   640
RB2  29   30   640
RB3  30   31   640
RB4  31   32   640
RB5  32   33   640
RB6  33   34   640
RB7  34   13   640
Q9   21   7    6    QN
Q10  22   29   6    QN
Q11  23   30   6    QN
Q12  24   31   6    QN
Q13  25   32   6    QN
Q14  26   33   6    QN
Q15  27   34   6    QN
Q16  28   13   6    QN
RC   40   41   15E6
CCTL 40   41   10.610E-15
I1   6    50   1.8E-3
R1   99   1    243.153
R2   99   4    243.153
*
* GAIN STAGE AND DOMINANT POLE AT 273HZ
*
EREF 98   0    POLY(2) (99,0) (50,0) 0 0.5 0.5
G1   98   8    (4,1) 4.113E-3
R5   8    98   243.153E6
C1   8    98   24E-13
V1   99   9    3.2
V2   10   50   3.2
D1   8    9    DX
D2   10   8    DX
*
* POLE AT 100MHZ
*
G5   98   35   (8,98) 1E-6
R11  35   98   1E6
C2   35   98   1.592E-15
*
* POLE AT 100MHZ
*
G6   98   36   (35,98) 1E-6
R12  36   98   1E6
C4   36   98   1.592E-15
*
* COMMON MODE GAIN STAGE WITH ZERO AT 200KHZ
*
ECM  37   98   (5,98) 1
R13  37   38   71.536
R14  38   98   1
C5   37   38   11.124E-9
*
* POLE AT 200MHZ
*
G3   98   45   (36,98) 1E-6
R10  45   98   1E6
C3   45   98   .796E-15
RGAT 70   98   30E3
MSW  45   71   98   50   MSWITCH
EGAT 71   98   POLY(1) (70,98) -5 3
*
* OUTPUT STAGE
*
GSY  99   50   POLY(1) (99,50) -11E-3 1.1E-3
FSY  99   50   POLY(2) V7 V8 21.2E-3 1 1
RO1  99   48   4
RO2  48   50   4
GO1  48   99   (99,45) 250E-3
GO2  50   48   (45,50) 250E-3
V4   48   46   -.516
V5   47   48   -.516
D5   46   45   DX
D6   45   47   DX
G4   98   44   (48,45) 250E-3
D7   44   42   DX
D8   43   44   DX
V7   42   98   0
V8   98   43   0
RF   11   48   2.242E3
RIN  11   2    20
.MODEL DX D(IS=1E-16)
.MODEL QN NPN(BF=1000)
.MODEL MSWITCH NMOS(VTO=2 W=100U L=10U KP=20)
.ENDS AD600J
