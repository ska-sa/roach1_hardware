* AD705T SPICE Macro-model 9/91, Rev. B
* AAG / PMI
*
* This version of the AD705 model simulates the worst case 
* parameters of the 'T' grade.  The worst case parameters
* used correspond to those in the data sheet.
*
* Revision History:
* REV B
* Updated op amp architecture
*
* Refer to "README.DOC" file for License Statement.  
* Use of this model indicates your acceptance with 
* the terms and provisions in the License Statement.
*
* Node assignments
*             non-inverting input
*             | inverting input
*             | |  positive supply
*             | |  |  negative supply
*             | |  |  |  output
*             | |  |  |  |  compensation
*             | |  |  |  |  |
.SUBCKT AD705T 1 2 99 50 31 15
*
* INPUT STAGE & POLE AT 3 MHz
*
IOS 1 2 DC 50E-12
CIN 1 2 2E-12
R1 2 3 2.586E8
R2 1 3 2.586E8
EOS 9 1 POLY(1) 19 25 25E-6 1
D1 2 9 DX
D2 9 2 DX
Q1 5 2 4 QX
Q2 6 9 4 QX
R3 99 5 1.5111E3
R4 99 6 1.5111E3
C2 5 6 17.554E-12
I1 4 50 34.227E-6
*
* FIRST GAIN STAGE
*
EREF 98 0 25 0 1
G1 98 12 5 6 57.46E-6
R7 12 98 1.4762E6
E1 99 13 POLY(1) 99 25 -2.4 1
D3 12 13 DX
E2 14 50 POLY(1) 25 50 -2.4 1
D4 14 12 DX
*
* SECOND GAIN STAGE & DOMINANT POLE AT 1.5 HZ
*
G2 98 15 12 25 11.409E-6
R8 15 98 310E6
C3 15 98 342.27E-12
V1 99 16 DC 2.3625
D5 15 16 DX
V2 17 50 DC 2.3625
D6 17 15 DX
*
* COMMON-MODE GAIN NETWORK WITH ZERO AT 4 kHz
*
ECM 18 98 3 25 1.9953
RCM1 18 19 1E6
CCM 18 19 39.88E-12
RCM2 19 98 1
*
* ZERO-POLE PAIR AT 165 kHz / 430 kHz
*
GZP 98 20 15 25 1E-6
RZP1 20 21 1E6
RZP2 21 98 1.6061E6
LZP 21 98 594.45E-3
*
* NEGATIVE ZERO AT -3 MHz
*
ENZ 22 98 20 25 1E6
RNZ1 22 23 1
CNZ 22 23 -53.052E-9
RNZ2 23 98 1E-6
*
* POLE AT 10 MHz
*
G3 98 24 23 25 1E-6
R9 24 98 1E6
C5 24 98 15.915E-15
*
* OUTPUT STAGE
*
IDC 99 50 DC 550.77E-6
RDC1 99 25 1E6
RDC2 25 50 1E6
DO1 99 26 DX
GO1 26 50 30 24 2E-3
DO2 50 26 DY
DO3 99 27 DX
GO2 27 50 24 30 2E-3
DO4 50 27 DY
VSC1 28 30 DC 3.15
DSC1 24 28 DX
VSC2 30 29 DC 3.15
DSC2 29 24 DX
GO3 30 99 99 24 2E-3
GO4 50 30 24 50 2E-3
RO1 99 30 500
RO2 30 50 500
LO 30 31 265E-9
*
* MODELS USED
*
.MODEL QX NPN(BF=1.7114E5)
.MODEL DX D(IS=1E-15)
.MODEL DY D(IS=1E-15 BV=50)
.ENDS AD705T
