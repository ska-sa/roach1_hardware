* OP481 SPICE Macro-model
* 7/97, Ver. 1
* TAM / ADSC
*
* Copyright 1996,1997 by Analog Devices
*
* Refer to "README.DOC" file for License Statement.  Use of this
* model indicates your acceptance of the terms and provisions in
* the License Statement.
*
* Node Assignments
*		noninverting input
*		|	inverting input
*		|	|	 positive supply
*		|	|	 |	 negative supply
*		|	|	 |	 |	 output
*		|	|	 |	 |	 |
*		|	|	 |	 |	 |
.SUBCKT OP481	1	2	99	50	45
*
* INPUT STAGE
*
Q1   4  1 3 PIX
Q2   6  7 5 PIX
I1  99  8 1.28E-6
EOS  7  2 POLY(1) (12,98) 80E-6 1
IOS  1  2 1E-10
RC1  4 50 500E3
RC2  6 50 500E3
RE1  3  8 108
RE2  5  8 108
V1  99 13 DC .9
V2  99 14 DC .9
D1   3 13 DX
D2   5 14 DX
*
* CMRR 76dB, ZERO AT 1kHz
*
ECM1 11 98 POLY(2) (1,98) (2,98) 0 .5 .5
R1   11 12 1.59E6
C1   11 12 100E-12
R2   12 98 283
*
* POLE AT 900kHz
*
EREF 98  0 (90,0) 1
G1   98 20 (4,6) 1E-6
R3   20 98 1E6
C2   20 98 177E-15
*
* POLE AT 500kHz
*
E2   21 98 (20,98) 1
R4   21 22 1E6
C3   22 98 320E-15
*
* GAIN STAGE
*
CF  45 40 8.5E-12
R5  40 98 65.65E6
G3  98 40 (22,98) 4.08E-7
D3  40 41 DX
D4  42 40 DX
V3  99 41 DC 0.5
V4  42 50 DC 0.5
*
* OUTPUT STAGE
*
ISY  99 50 1.375E-6
RS1  99 90 10E6
RS2  90 50 10E6
M1  48 46 99 99 POX L=1.5u W=300u
M2  49 47 50 50 NOX L=1.5u W=300u
RO1 48 45 400
RO2 49 45 200
EG1 99 46 POLY(1) (98,40) 0.77 1
EG2 47 50 POLY(1) (40,98) 0.77 1
*
* MODELS
*
.MODEL POX PMOS (LEVEL=2, KP=25E-6, VTO=-0.75, LAMBDA=0.01)
.MODEL NOX NMOS (LEVEL=2, KP=25E-6, VTO=0.75,  LAMBDA=0.01)
.MODEL PIX PNP (BF=200)
.MODEL DX D(IS=1E-14)
.ENDS OP481