* AD829S SPICE Macro-model                   9/90, Rev. A
*                                            JCB / PMI
*
* This version of the AD829 model simulates the worst case 
* parameters of the 'S' grade.  The worst case parameters
* used correspond to those in the data sheet.
*
* Copyright 1990 by Analog Devices
*
* Refer to "README.DOC" file for License Statement.  Use of this model
* indicates your acceptance with the terms and provisions in the License Statement.
*
* Node assignments
*               non-inverting input
*               | inverting input
*               | | positive supply
*               | | |  negative supply
*               | | |  |  output
*               | | |  |  |  compensation node
*               | | |  |  |  |
.SUBCKT AD829S  1 2 99 50 30 12
*
* INPUT STAGE & POLE AT 200 MHZ
*
R1   2  3     17.8E3
R2   1  3     17.8E3
R3   5 99     56.4
R4   6 99     56.4
CIN  1  2     5E-12
C2   5  6     7.18E-12
I1   4  50    1.2E-3
IOS  1  2     250E-9
EOS  9  1     POLY(1)  19 23  0.5E-3  1
Q1   5  2 10  QX
Q2   6  9 11  QX
R5   10 4     13.4
R6   11 4     13.4
*
EREF 98 0     23  0  1
*
* GAIN STAGE & DOMINANT POLE AT 2.7 KHZ
*
R7  12 98     2.82E6
C3  12 98     5.2E-12
G1  98 12     5  6  17.73E-3
V2  99 13     3.4
V3  14 50     3.4
D3  12 13     DX
D4  14 12     DX
*
* ZERO/POLE PAIR AT 50MHz/100MHz
*
R8  15 16     1E6
R9  16 98     1E6
L1  16 98     1.59E-3
G2  98 15     12 23  1E-6
*
* POLE AT 400 MHZ
*
R41 41 98     1E6
C41 41 98     398E-18
G41 98 41     15 23  1E-6
*
* POLE AT 400 MHZ
*
R42 42 98     1E6
C42 42 98     398E-18
G42 98 42     41 23  1E-6
*
* POLE AT 200 MHZ
*
R43 43 98     1E6
C43 43 98     796E-18
G43 98 43     42 23  1E-6
*
* COMMON-MODE GAIN NETWORK WITH ZERO AT 30 KHZ
*
R11 18 19     1E6
C6  18 19     5.31E-12
R12 19 98     1
E2  18 98     3  23  10
*
* POLE AT 400 MHZ
*
R15 22 98     1E6
C8  22 98     398E-18
G3  98 22     43 23  1E-6
*
* OUTPUT STAGE
*
RF  25 60     500
CF  60 12     12.5E-12
R16 23 99     100E3
R17 23 50     100E3
ISY 99 50     5.45E-3
R18 25 99     30
R19 25 50     30
L2  25 30     1E-8
G4  28 50     22 25  33.33E-3
G5  29 50     25 22  33.33E-3
G6  25 99     99 22  33.33E-3
G7  50 25     22 50  33.33E-3
V4  26 25     -0.2
V5  25 27     -0.2
D5  22 26     DX
D6  27 22     DX
D7  99 28     DX
D8  99 29     DX
D9  50 28     DY
D10 50 29     DY
*
* MODELS USED
*
.MODEL QX NPN(BF=85.7)
.MODEL DX   D(IS=1E-15)
.MODEL DY   D(IS=1E-15 BV=50)
.ENDS
