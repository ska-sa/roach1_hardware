**/////////////////////////////////////////////////////////////////////////////
**$Date: 2007/11/06 18:10:54 $
**$RCSfile: v5_gtp_voltage_settings_slow.ckt,v $
**$Revision: 1.1 $
**//////////////////////////////////////////////////////////////////////////////
**   ____  ____ 
**  /   /\/   / 
** /___/  \  /    Vendor: Xilinx 
** \   \   \/     Version : 1.0
**  \   \         Filename : v5_gtp_voltage_settings_slow.ckt
**  /   /         
** /___/   /\
** \   \  /  \ 
**  \___\/\___\ 
**
**                VIRTEX-5 FPGA ROCKETIO SIGNAL INTEGRITY KIT
**
**
** Description : Virtex-5 GTP Transmit and Receive Analog and Threshold 
**               Supply Voltage Settings for slow operating conditions
**//////////////////////////////////////////////////////////////////////////////

** Virtex-5 GTP Transmitter Voltages **
.param vsup_tx_v5_gtp  = 0.95
.param vsuph_tx_v5_gtp = 1.14

** Virtex-5 GTP Receiver Voltages **
.param vsup_rx_v5_gtp  = 0.95
.param vsuph_rx_v5_gtp = 1.14

** Virtex-5 GTP Refclk Voltages **
.param vsup_refclk_v5_gtp  = 0.95
.param vsuph_refclk_v5_gtp = 1.14