* Netlist for net Lsw00 - D:\ROACH\elec\SISim\roach_ddr2_dqs_single_fpga2dimm.sp


* Output from HyperLynx SPICE Writer
* Created by Francois on Date: Wednesday Nov. 28,2007   Time: 15:33:06
* Created with HyperLynx version: 7.7 build: 385
* Design file: roach_ddr2_dq_dual_fpga2dimm.ffs
* Special Settings: Coupled


.SUBCKT roach_ddr2_dqs_single_fpga2dimm Vinp Vinn 100 105 131 107 111 132 115 133 119 134 126 135 128 136

* Node  #  = <Reference Designator>.<pin name>
**********************************************
* Node 100 = J1.Port4 (at pin)
* Node 105 = U8.1 (at pin) (receiver)
X_mdl_105 105 d_receive_105 MODEL_U8_1_ip
* Node 131 = R8.1 (at pin)
* Node 107 = J1.Port3 (at pin)
* Node 111 = R7.2 (at pin)
* Node 132 = U7.1 (at pin) (receiver)
X_mdl_113 113 d_receive_113 MODEL_U7_1_ip
* Node 115 = J1.Port2 (at pin)
* Node 133 = U6.1 (at pin) (driver)
X_mdl_117 117 Vinn MODEL_U6_1_ip
* Node 119 = J1.Port1 (at pin)
* Node 134 = U5.1 (at pin) (driver)
X_mdl_121 121 Vinp MODEL_U5_1_ip
* Node 126 = U3.2 (at pin) (driver)
X_mdl_124 124 Vinn MODEL_U3_2_ip
* Node 135 = R1.2 (at pin)
* Node 128 = R1.1 (at pin)
* Node 136 = U3.1 (at pin) (driver)
X_mdl_129 129 Vinp MODEL_U3_1_ip

* Node   0 = Gnd (Common Return)

.connect 136 128 

.connect 135 126 

.connect 134 119 

.connect 133 115 

.connect 132 111 

.connect 131 105 


CV001       102    0 3.645e-013
R8_1        105    4 50
CV002       109    0 3.645e-013
TP012       111    0  113    0 Z0=1.171893e+002 TD=1.757840e-011
R7_2        111    4 50
TP013       115    0  117    0 Z0=3.579990e+001 TD=8.770975e-011
TP014       119    0  121    0 Z0=3.579990e+001 TD=8.770975e-011
TP015       126    0  124    0 Z0=3.579990e+001 TD=8.770975e-011
R1_2        126  128 50
TP018       128    0  129    0 Z0=3.579990e+001 TD=8.770975e-011

WCond_000  102 109 0 105 111 0 RLGCmodel=Cond_000 N=2 L=0.050000 fgd=1e9  MULTIDEBYE=1
WCond_001  107 100 0 109 102 0 RLGCmodel=Cond_001 N=2 L=0.005000 fgd=1e9  MULTIDEBYE=1
V4  4  0  0.90
V3  3  0  1.00
V2  2  0  1.80
V1  1  0  0.00

****  Transmission line models ***********************
*********************************
* RLGC model created by HyperLynx SPICE generator
*
.MODEL Cond_000 W MODELTYPE=RLGC N=2
* Lo  (H/m)
+ Lo =
+ 5.18283e-007  
+ 1.07974e-007  5.18283e-007  

* Co  (F/m)
+ Co =
+ 9.65006e-011  
+ -2.01039e-011  9.65006e-011  

* Loss turned off.  Only lossless components written.

*********************************

*********************************
* RLGC model created by HyperLynx SPICE generator
*
.MODEL Cond_001 W MODELTYPE=RLGC N=2
* Lo  (H/m)
+ Lo =
+ 5.50676e-007  
+ 2.16403e-007  5.50676e-007  

* Co  (F/m)
+ Co =
+ 6.99599e-011  
+ -2.34655e-011  6.99599e-011  

* Loss turned off.  Only lossless components written.

*********************************

****  End Transmission line models *******************

.ENDS

* IBIS model subcircuit definitions
**********************************************
*Define subcircuit for MODEL_U8_1_ip
.subckt MODEL_U8_1_ip a_signal d_receive 
VPullUpRef a_PURef 0 1.8
VPullDownRef a_PDRef 0 0

X_105 a_signal d_receive 0 a_PURef a_PDRef MODEL_U8_1

.ends MODEL_U8_1_ip

*Define subcircuit for MODEL_U8_1
.subckt MODEL_U8_1 a_signal d_receive a_gnd a_PURef a_PDRef 

C_comp a_signal a_gnd 2.811e-012

VGCRef a_GCRef 0 0
G_gnd_clamp a_signal a_GCRef table v(a_signal, a_GCRef) = 
+ (-23.4,-22.2654) (-1.8,-0.760219) (-1.795,-0.755241) 
+ (-1.79,-0.750299) (-1.785,-0.745359) (-1.78,-0.740421) 
+ (-1.775,-0.735484) (-1.77,-0.730549) (-1.765,-0.725617) 
+ (-1.755,-0.715754) (-1.735,-0.696055) (-1.73,-0.691139) 
+ (-1.695,-0.656751) (-1.69,-0.651848) (-1.63,-0.593191) 
+ (-1.625,-0.588303) (-1.62,-0.583444) (-1.615,-0.578597) 
+ (-1.55,-0.51558) (-1.545,-0.510732) (-1.54,-0.505913) 
+ (-1.53,-0.496355) (-1.525,-0.491576) (-1.45,-0.419894) 
+ (-1.445,-0.415115) (-1.44,-0.410336) (-1.435,-0.40558) 
+ (-1.415,-0.387037) (-1.41,-0.382402) (-1.32,-0.29896) 
+ (-1.315,-0.294325) (-1.3,-0.280418) (-1.295,-0.275794) 
+ (-1.27,-0.254226) (-1.265,-0.249912) (-1.175,-0.172264) 
+ (-1.17,-0.16795) (-1.16,-0.159323) (-1.155,-0.155515) 
+ (-1.14,-0.145365) (-1.135,-0.141982) (-1.04,-0.0776975) 
+ (-1.035,-0.0743141) (-1.01,-0.0573972) (-1.005,-0.0557414) 
+ (-0.98,-0.0484965) (-0.975,-0.0470476) (-0.94,-0.0369047) 
+ (-0.935,-0.0354557) (-0.895,-0.0238639) (-0.89,-0.0230547) 
+ (-0.875,-0.0215177) (-0.87,-0.0210053) (-0.825,-0.0163943) 
+ (-0.82,-0.0158819) (-0.795,-0.0133202) (-0.79,-0.0128917) 
+ (-0.78,-0.0122114) (-0.775,-0.0118712) (-0.745,-0.00983015) 
+ (-0.74,-0.00948997) (-0.7,-0.00676859) (-0.695,-0.0065163) 
+ (-0.69,-0.00628185) (-0.685,-0.0060474) (-0.65,-0.00440625) 
+ (-0.645,-0.00417181) (-0.615,-0.00276511) (-0.61,-0.00255864) 
+ (-0.605,-0.0024436) (-0.56,-0.00140824) (-0.555,-0.0012932) 
+ (-0.535,-0.000833048) (-0.53,-0.000718009) (-0.525,-0.00064001) 
+ (-0.515,-0.000581028) (-0.51,-0.000551537) (-0.49,-0.000433574) 
+ (-0.485,-0.000404083) (-0.475,-0.000345101) (-0.47,-0.00031561) 
+ (-0.44,-0.000138664) (-0.435,-0.000122592) (-0.41,-9.27216e-005) 
+ (-0.39,-6.88249e-005) (-0.385,-6.50985e-005) (-0.365,-5.80787e-005) 
+ (-0.355,-5.45688e-005) (-0.35,-5.28139e-005) (-0.325,-4.40391e-005) 
+ (-0.32,-4.25496e-005) (-0.285,0) (3.6,0) 
+ (25.2,0) 

VPCRef a_PCRef 0 1.8
G_power_clamp a_PCRef a_signal table v(a_PCRef, a_signal) = 
+ (-23.4,-18.3) (-1.8,-0.607667) (-1.795,-0.603572) 
+ (-1.79,-0.599504) (-1.785,-0.595438) (-1.78,-0.591374) 
+ (-1.775,-0.587311) (-1.77,-0.58325) (-1.765,-0.57919) 
+ (-1.755,-0.571074) (-1.735,-0.554862) (-1.73,-0.550816) 
+ (-1.695,-0.522518) (-1.69,-0.518485) (-1.63,-0.470223) 
+ (-1.625,-0.466201) (-1.62,-0.462204) (-1.615,-0.458217) 
+ (-1.55,-0.406381) (-1.545,-0.402394) (-1.54,-0.39843) 
+ (-1.53,-0.390572) (-1.525,-0.386643) (-1.45,-0.327709) 
+ (-1.445,-0.32378) (-1.44,-0.319851) (-1.435,-0.315941) 
+ (-1.415,-0.300718) (-1.41,-0.296913) (-1.32,-0.228411) 
+ (-1.315,-0.224606) (-1.3,-0.213189) (-1.295,-0.209394) 
+ (-1.27,-0.191808) (-1.265,-0.188291) (-1.175,-0.124981) 
+ (-1.17,-0.121464) (-1.16,-0.114429) (-1.155,-0.111406) 
+ (-1.14,-0.103581) (-1.135,-0.100972) (-1.04,-0.0514083) 
+ (-1.035,-0.0487997) (-1.01,-0.0357566) (-1.005,-0.0346027) 
+ (-0.98,-0.0297033) (-0.975,-0.0287235) (-0.94,-0.0218644) 
+ (-0.935,-0.0208845) (-0.895,-0.0130456) (-0.89,-0.0124844) 
+ (-0.875,-0.0113837) (-0.87,-0.0110168) (-0.825,-0.0077146) 
+ (-0.82,-0.0073477) (-0.795,-0.00551317) (-0.79,-0.00523633) 
+ (-0.78,-0.00487255) (-0.775,-0.00469066) (-0.745,-0.00359931) 
+ (-0.74,-0.00341742) (-0.7,-0.0019623) (-0.695,-0.00186186) 
+ (-0.69,-0.00177795) (-0.685,-0.00169404) (-0.65,-0.00110668) 
+ (-0.645,-0.00102277) (-0.615,-0.000519312) (-0.61,-0.000449671) 
+ (-0.605,-0.000426662) (-0.56,-0.000219585) (-0.555,-0.000196577) 
+ (-0.535,-0.000104543) (-0.53,-8.15342e-005) (-0.525,-6.69439e-005) 
+ (-0.515,-5.98123e-005) (-0.51,-5.62465e-005) (-0.49,-4.19832e-005) 
+ (-0.475,-3.12858e-005) (-0.47,-2.77199e-005) (-0.44,-6.32505e-006) 
+ (-0.435,-4.48769e-006) (-0.41,-1.80397e-006) (-0.393,0) 
+ (3.6,0) (25.2,0) 

* IBIS style receiver logic.  No hysteresis.
Y_rx_logic ibis_receiver_logic(icx_behavioral)
+ GENERIC: corner="ibis_typ"
+          vinL_values="(0.650000,0.650000,0.650000)"
+          vinH_values="(1.150000,1.150000,1.150000)"
+ PORT: a_gnd
+       a_signal
+       d_receive

.model ibis_receiver_logic(icx_behavioral) MACRO LANG=VHDLAMS LIB=icxbase
.ends MODEL_U8_1

*Define subcircuit for MODEL_U7_1_ip
.subckt MODEL_U7_1_ip a_signal d_receive 
VPullUpRef a_PURef 0 1.8
VPullDownRef a_PDRef 0 0

X_132 a_signal d_receive 0 a_PURef a_PDRef MODEL_U7_1

.ends MODEL_U7_1_ip

*Define subcircuit for MODEL_U7_1
.subckt MODEL_U7_1 a_signal d_receive a_gnd a_PURef a_PDRef 

C_comp a_signal a_gnd 2.811e-012

VGCRef a_GCRef 0 0
G_gnd_clamp a_signal a_GCRef table v(a_signal, a_GCRef) = 
+ (-23.4,-22.2654) (-1.8,-0.760219) (-1.795,-0.755241) 
+ (-1.79,-0.750299) (-1.785,-0.745359) (-1.78,-0.740421) 
+ (-1.775,-0.735484) (-1.77,-0.730549) (-1.765,-0.725617) 
+ (-1.755,-0.715754) (-1.735,-0.696055) (-1.73,-0.691139) 
+ (-1.695,-0.656751) (-1.69,-0.651848) (-1.63,-0.593191) 
+ (-1.625,-0.588303) (-1.62,-0.583444) (-1.615,-0.578597) 
+ (-1.55,-0.51558) (-1.545,-0.510732) (-1.54,-0.505913) 
+ (-1.53,-0.496355) (-1.525,-0.491576) (-1.45,-0.419894) 
+ (-1.445,-0.415115) (-1.44,-0.410336) (-1.435,-0.40558) 
+ (-1.415,-0.387037) (-1.41,-0.382402) (-1.32,-0.29896) 
+ (-1.315,-0.294325) (-1.3,-0.280418) (-1.295,-0.275794) 
+ (-1.27,-0.254226) (-1.265,-0.249912) (-1.175,-0.172264) 
+ (-1.17,-0.16795) (-1.16,-0.159323) (-1.155,-0.155515) 
+ (-1.14,-0.145365) (-1.135,-0.141982) (-1.04,-0.0776975) 
+ (-1.035,-0.0743141) (-1.01,-0.0573972) (-1.005,-0.0557414) 
+ (-0.98,-0.0484965) (-0.975,-0.0470476) (-0.94,-0.0369047) 
+ (-0.935,-0.0354557) (-0.895,-0.0238639) (-0.89,-0.0230547) 
+ (-0.875,-0.0215177) (-0.87,-0.0210053) (-0.825,-0.0163943) 
+ (-0.82,-0.0158819) (-0.795,-0.0133202) (-0.79,-0.0128917) 
+ (-0.78,-0.0122114) (-0.775,-0.0118712) (-0.745,-0.00983015) 
+ (-0.74,-0.00948997) (-0.7,-0.00676859) (-0.695,-0.0065163) 
+ (-0.69,-0.00628185) (-0.685,-0.0060474) (-0.65,-0.00440625) 
+ (-0.645,-0.00417181) (-0.615,-0.00276511) (-0.61,-0.00255864) 
+ (-0.605,-0.0024436) (-0.56,-0.00140824) (-0.555,-0.0012932) 
+ (-0.535,-0.000833048) (-0.53,-0.000718009) (-0.525,-0.00064001) 
+ (-0.515,-0.000581028) (-0.51,-0.000551537) (-0.49,-0.000433574) 
+ (-0.485,-0.000404083) (-0.475,-0.000345101) (-0.47,-0.00031561) 
+ (-0.44,-0.000138664) (-0.435,-0.000122592) (-0.41,-9.27216e-005) 
+ (-0.39,-6.88249e-005) (-0.385,-6.50985e-005) (-0.365,-5.80787e-005) 
+ (-0.355,-5.45688e-005) (-0.35,-5.28139e-005) (-0.325,-4.40391e-005) 
+ (-0.32,-4.25496e-005) (-0.285,0) (3.6,0) 
+ (25.2,0) 

VPCRef a_PCRef 0 1.8
G_power_clamp a_PCRef a_signal table v(a_PCRef, a_signal) = 
+ (-23.4,-18.3) (-1.8,-0.607667) (-1.795,-0.603572) 
+ (-1.79,-0.599504) (-1.785,-0.595438) (-1.78,-0.591374) 
+ (-1.775,-0.587311) (-1.77,-0.58325) (-1.765,-0.57919) 
+ (-1.755,-0.571074) (-1.735,-0.554862) (-1.73,-0.550816) 
+ (-1.695,-0.522518) (-1.69,-0.518485) (-1.63,-0.470223) 
+ (-1.625,-0.466201) (-1.62,-0.462204) (-1.615,-0.458217) 
+ (-1.55,-0.406381) (-1.545,-0.402394) (-1.54,-0.39843) 
+ (-1.53,-0.390572) (-1.525,-0.386643) (-1.45,-0.327709) 
+ (-1.445,-0.32378) (-1.44,-0.319851) (-1.435,-0.315941) 
+ (-1.415,-0.300718) (-1.41,-0.296913) (-1.32,-0.228411) 
+ (-1.315,-0.224606) (-1.3,-0.213189) (-1.295,-0.209394) 
+ (-1.27,-0.191808) (-1.265,-0.188291) (-1.175,-0.124981) 
+ (-1.17,-0.121464) (-1.16,-0.114429) (-1.155,-0.111406) 
+ (-1.14,-0.103581) (-1.135,-0.100972) (-1.04,-0.0514083) 
+ (-1.035,-0.0487997) (-1.01,-0.0357566) (-1.005,-0.0346027) 
+ (-0.98,-0.0297033) (-0.975,-0.0287235) (-0.94,-0.0218644) 
+ (-0.935,-0.0208845) (-0.895,-0.0130456) (-0.89,-0.0124844) 
+ (-0.875,-0.0113837) (-0.87,-0.0110168) (-0.825,-0.0077146) 
+ (-0.82,-0.0073477) (-0.795,-0.00551317) (-0.79,-0.00523633) 
+ (-0.78,-0.00487255) (-0.775,-0.00469066) (-0.745,-0.00359931) 
+ (-0.74,-0.00341742) (-0.7,-0.0019623) (-0.695,-0.00186186) 
+ (-0.69,-0.00177795) (-0.685,-0.00169404) (-0.65,-0.00110668) 
+ (-0.645,-0.00102277) (-0.615,-0.000519312) (-0.61,-0.000449671) 
+ (-0.605,-0.000426662) (-0.56,-0.000219585) (-0.555,-0.000196577) 
+ (-0.535,-0.000104543) (-0.53,-8.15342e-005) (-0.525,-6.69439e-005) 
+ (-0.515,-5.98123e-005) (-0.51,-5.62465e-005) (-0.49,-4.19832e-005) 
+ (-0.475,-3.12858e-005) (-0.47,-2.77199e-005) (-0.44,-6.32505e-006) 
+ (-0.435,-4.48769e-006) (-0.41,-1.80397e-006) (-0.393,0) 
+ (3.6,0) (25.2,0) 

* IBIS style receiver logic.  No hysteresis.
Y_rx_logic ibis_receiver_logic(icx_behavioral)
+ GENERIC: corner="ibis_typ"
+          vinL_values="(0.650000,0.650000,0.650000)"
+          vinH_values="(1.150000,1.150000,1.150000)"
+ PORT: a_gnd
+       a_signal
+       d_receive

.model ibis_receiver_logic(icx_behavioral) MACRO LANG=VHDLAMS LIB=icxbase
.ends MODEL_U7_1

*Define subcircuit for MODEL_U6_1_ip
.subckt MODEL_U6_1_ip a_signal a_control 
VPullUpRef a_PURef 0 1.8
VPullDownRef a_PDRef 0 1e-100


Y_a_control ibis_driver_logic(icx_behavioral)
+ GENERIC: corner="ibis_typ"
+          vmeas_values="( 0.5, 0.5, 0.5 )"
+ PORT: a_control
+       a_gnd
+       d_control

.model ibis_driver_logic(icx_behavioral) MACRO LANG=VHDLAMS LIB=icxbase

X_133 a_signal d_control 0 a_PURef a_PDRef MODEL_U6_1

.ends MODEL_U6_1_ip

*Define subcircuit for MODEL_U6_1
.subckt MODEL_U6_1 a_signal d_control a_gnd a_PURef a_PDRef

C_comp a_signal a_gnd 6e-012

VGCRef a_GCRef 0 0
G_gnd_clamp a_signal a_GCRef table v(a_signal, a_GCRef) = 
+ (-3,0) (1,0) (2,0) 
+ (6,0) 

VPCRef a_PCRef 0 1.8
G_power_clamp a_PCRef a_signal table v(a_PCRef, a_signal) = 
+ (-6,0) (-2,0) (-1,0) 
+ (3,0) 

Y_control ibis_control(icx_behavioral)
+ PORT: d_control
+       d_pullup_control
+       d_pulldown_control

.model ibis_control(icx_behavioral) MACRO LANG=VHDLAMS LIB=icxbase


*IBIS Pulldown tables
Y_PullDown ibis_ktiv(icx_behavioral)
+ GENERIC: corner="ibis_typ"
+          tdata_0to1_typ="(1.63161e-011, 2.2246e-011, 2.81759e-011, 3.41058e-011, 4.00356e-011, 4.59655e-011,
+ 5.18954e-011, 5.78253e-011, 6.37551e-011, 6.9685e-011, 7.56149e-011, 8.15448e-011,
+ 8.74746e-011, 9.34045e-011, 9.93344e-011, 1.05264e-010, 1.11194e-010, 1.17124e-010,
+ 1.23054e-010, 1.28984e-010, 1.34914e-010, 1.40843e-010, 1.46773e-010, 1.52703e-010,
+ 1.58633e-010, 1.64563e-010, 1.70493e-010, 1.76423e-010, 1.82353e-010, 1.88282e-010,
+ 1.94212e-010, 2.00142e-010, 2.06072e-010, 2.12002e-010, 2.17932e-010, 2.23862e-010,
+ 2.29792e-010, 2.35721e-010, 2.41651e-010, 2.47581e-010, 2.53511e-010, 2.59441e-010,
+ 2.65371e-010, 2.71301e-010, 2.77231e-010, 2.8316e-010, 2.8909e-010, 2.9502e-010,
+ 3.0095e-010, 3.0688e-010, 3.1281e-010, 3.1874e-010, 3.2467e-010, 3.30599e-010,
+ 3.36529e-010, 3.42459e-010, 3.48389e-010, 3.54319e-010, 3.60249e-010, 3.66179e-010,
+ 3.72109e-010, 3.78038e-010, 3.83968e-010, 3.89898e-010, 3.95828e-010, 4.01758e-010,
+ 4.07688e-010, 4.13618e-010, 4.19548e-010, 4.25477e-010, 4.31407e-010, 4.37337e-010,
+ 4.43267e-010, 4.49197e-010, 4.55127e-010, 4.61057e-010, 4.66987e-010, 4.72916e-010,
+ 4.78846e-010, 4.84776e-010, 4.90706e-010, 4.96636e-010, 5.02566e-010, 5.08496e-010,
+ 5.14426e-010, 5.20355e-010, 5.26285e-010, 5.32215e-010, 5.38145e-010, 5.44075e-010,
+ 5.50005e-010, 5.55935e-010, 5.61865e-010, 5.67794e-010, 5.73724e-010, 5.79654e-010,
+ 5.85584e-010, 5.91514e-010, 5.97444e-010, 6.03374e-010, 6.09304e-010, 6.15233e-010,
+ 6.21163e-010, 6.27093e-010, 6.33023e-010, 6.38953e-010, 6.44883e-010, 6.50813e-010,
+ 6.56743e-010, 6.62672e-010, 6.68602e-010, 6.74532e-010, 6.80462e-010, 6.86392e-010,
+ 6.92322e-010, 6.98252e-010, 7.04182e-010, 7.10111e-010, 7.16041e-010, 7.21971e-010,
+ 7.27901e-010, 7.33831e-010, 7.39761e-010, 7.45691e-010, 7.51621e-010, 7.5755e-010,
+ 7.6348e-010, 7.6941e-010, 7.7534e-010, 7.8127e-010, 7.872e-010, 7.9313e-010,
+ 7.9906e-010, 8.04989e-010, 8.10919e-010, 8.16849e-010, 8.22779e-010, 8.28709e-010,
+ 8.34639e-010, 8.40569e-010, 8.46499e-010, 8.52428e-010, 8.58358e-010, 8.64288e-010,
+ 8.70218e-010, 8.76148e-010, 8.82078e-010, 8.88008e-010, 8.93938e-010, 8.99867e-010,
+ 9.05797e-010, 9.11727e-010, 9.17657e-010, 9.23587e-010, 9.29517e-010, 9.35447e-010,
+ 9.41377e-010, 9.47306e-010, 9.53236e-010, 9.59166e-010, 9.65096e-010, 9.71026e-010,
+ 9.76956e-010, 9.82886e-010, 9.88816e-010, 9.94745e-010, 1.00068e-009, 1.00661e-009,
+ 1.01254e-009, 1.01846e-009, 1.02439e-009, 1.03032e-009, 1.03625e-009, 1.04218e-009,
+ 1.04811e-009, 1.05404e-009, 1.05997e-009, 1.0659e-009, 1.07183e-009, 1.07776e-009,
+ 1.08369e-009, 1.08962e-009, 1.09555e-009, 1.10148e-009, 1.10741e-009, 1.11334e-009,
+ 1.11927e-009, 1.1252e-009, 1.13113e-009, 1.13706e-009, 1.14299e-009, 1.14892e-009,
+ 1.15485e-009, 1.16078e-009, 1.16671e-009, 1.17264e-009, 1.17857e-009, 1.1845e-009,
+ 1.19043e-009, 1.19636e-009, 1.20229e-009, 1.20822e-009)"
+          kdata_0to1_typ="(0, 0.00693597, 0.00734267, 0.00775038, 0.00815913, 0.00858505,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0.0149774, 0.0168403, 0.0186985, 0.0205519,
+ 0.0224006, 0.0240851, 0.0257124, 0.0534193, 0.0575498, 0.0616171,
+ 0.0656214, 0.069563, 0.102944, 0.109289, 0.1155, 0.121575,
+ 0.127512, 0.185885, 0.194014, 0.201885, 0.209487, 0.216904,
+ 0.262763, 0.270595, 0.278029, 0.284935, 0.291331, 0.389536,
+ 0.397239, 0.403807, 0.409531, 0.41272, 0.458302, 0.460574,
+ 0.460332, 0.45866, 0.456168, 0.521521, 0.519402, 0.516554,
+ 0.512182, 0.507981, 0.562714, 0.560143, 0.557616, 0.556013,
+ 0.55331, 0.659015, 0.662791, 0.666581, 0.669294, 0.672524,
+ 0.716442, 0.724711, 0.731962, 0.740509, 0.749691, 0.739752,
+ 0.749267, 0.759439, 0.770012, 0.780565, 0.791097, 0.79587,
+ 0.809271, 0.822809, 0.836161, 0.849325, 0.834494, 0.847778,
+ 0.862015, 0.876457, 0.891109, 0.864523, 0.877546, 0.890758,
+ 0.904235, 0.918949, 0.917735, 0.932302, 0.946993, 0.961955,
+ 0.977195, 0.924242, 0.935102, 0.946108, 0.957264, 0.968572,
+ 0.909004, 0.915836, 0.922722, 0.929662, 0.936656, 0.952113,
+ 0.960445, 0.968871, 0.977393, 0.986011, 0.960073, 0.966314,
+ 0.972606, 0.97895, 0.985348, 0.970999, 0.976042, 0.98112,
+ 0.986232, 0.991379, 0.972387, 0.975803, 0.979234, 0.98268,
+ 0.986141, 0.967094, 0.968918, 0.970746, 0.972578, 0.974414,
+ 0.973267, 0.97489, 0.976515, 0.978144, 0.979776, 0.98008,
+ 0.981606, 0.983135, 0.984771, 0.986428, 0.984285, 0.985785,
+ 0.987287, 0.988793, 0.990302, 0.982654, 0.983469, 0.984284,
+ 0.9851, 0.985918, 0.989565, 0.990614, 0.991664, 0.992715,
+ 0.993768, 0.993327, 0.994265, 0.995205, 0.996146, 0.997089,
+ 0.998032, 1, 1, 1, 1, 1,
+ 0.99667, 0.997028, 0.997387, 0.997745, 0.998104, 0.993811,
+ 0.993821, 0.99383, 0.99384, 0.993849, 0.998489, 0.998848,
+ 0.999207, 0.999566, 0.999926, 0.998882, 0.999149, 0.999417,
+ 0.999684, 0.999951, 1, 1)"
+          tdata_1to0_typ="(7.19709e-011, 7.82209e-011, 8.44709e-011, 9.07209e-011, 9.69709e-011, 1.03221e-010,
+ 1.09471e-010, 1.15721e-010, 1.21971e-010, 1.28221e-010, 1.34471e-010, 1.40721e-010,
+ 1.46971e-010, 1.53221e-010, 1.59471e-010, 1.65721e-010, 1.71971e-010, 1.78221e-010,
+ 1.84471e-010, 1.90721e-010, 1.96971e-010, 2.03221e-010, 2.09471e-010, 2.15721e-010,
+ 2.21971e-010, 2.28221e-010, 2.34471e-010, 2.40721e-010, 2.46971e-010, 2.53221e-010,
+ 2.59471e-010, 2.65721e-010, 2.71971e-010, 2.78221e-010, 2.84471e-010, 2.90721e-010,
+ 2.96971e-010, 3.03221e-010, 3.09471e-010, 3.15721e-010, 3.21971e-010, 3.28221e-010,
+ 3.34471e-010, 3.40721e-010, 3.46971e-010, 3.53221e-010, 3.59471e-010, 3.65721e-010,
+ 3.71971e-010, 3.78221e-010, 3.84471e-010, 3.90721e-010, 3.96971e-010, 4.03221e-010,
+ 4.09471e-010, 4.15721e-010, 4.21971e-010, 4.28221e-010, 4.34471e-010, 4.40721e-010,
+ 4.46971e-010, 4.53221e-010, 4.59471e-010, 4.65721e-010, 4.71971e-010, 4.78221e-010,
+ 4.84471e-010, 4.90721e-010, 4.96971e-010, 5.03221e-010, 5.09471e-010, 5.15721e-010,
+ 5.21971e-010, 5.28221e-010, 5.34471e-010, 5.40721e-010, 5.46971e-010, 5.53221e-010,
+ 5.59471e-010, 5.65721e-010, 5.71971e-010, 5.78221e-010, 5.84471e-010, 5.90721e-010,
+ 5.96971e-010, 6.03221e-010, 6.09471e-010, 6.15721e-010, 6.21971e-010, 6.28221e-010,
+ 6.34471e-010, 6.40721e-010, 6.46971e-010, 6.53221e-010, 6.59471e-010, 6.65721e-010,
+ 6.71971e-010, 6.78221e-010, 6.84471e-010, 6.90721e-010, 6.96971e-010, 7.03221e-010,
+ 7.09471e-010, 7.15721e-010, 7.21971e-010, 7.28221e-010, 7.34471e-010, 7.40721e-010,
+ 7.46971e-010, 7.53221e-010, 7.59471e-010, 7.65721e-010, 7.71971e-010, 7.78221e-010,
+ 7.84471e-010, 7.90721e-010, 7.96971e-010, 8.03221e-010, 8.09471e-010, 8.15721e-010,
+ 8.21971e-010, 8.28221e-010, 8.34471e-010, 8.40721e-010, 8.46971e-010, 8.53221e-010,
+ 8.59471e-010, 8.65721e-010, 8.71971e-010, 8.78221e-010, 8.84471e-010, 8.90721e-010,
+ 8.96971e-010, 9.03221e-010, 9.09471e-010, 9.15721e-010, 9.21971e-010, 9.28221e-010,
+ 9.34471e-010, 9.40721e-010, 9.46971e-010, 9.53221e-010, 9.59471e-010, 9.65721e-010,
+ 9.71971e-010, 9.78221e-010, 9.84471e-010, 9.90721e-010, 9.96971e-010, 1.00322e-009,
+ 1.00947e-009, 1.01572e-009, 1.02197e-009, 1.02822e-009, 1.03447e-009, 1.04072e-009,
+ 1.04697e-009, 1.05322e-009, 1.05947e-009, 1.06572e-009, 1.07197e-009, 1.07822e-009,
+ 1.08447e-009, 1.09072e-009, 1.09697e-009, 1.10322e-009, 1.10947e-009, 1.11572e-009,
+ 1.12197e-009, 1.12822e-009, 1.13447e-009, 1.14072e-009, 1.14697e-009, 1.15322e-009,
+ 1.15947e-009, 1.16572e-009, 1.17197e-009, 1.17822e-009, 1.18447e-009, 1.19072e-009,
+ 1.19697e-009, 1.20322e-009, 1.20947e-009, 1.21572e-009, 1.22197e-009, 1.22822e-009,
+ 1.23447e-009, 1.24072e-009, 1.24697e-009, 1.25322e-009, 1.25947e-009, 1.26572e-009,
+ 1.27197e-009, 1.27822e-009, 1.28447e-009, 1.29072e-009, 1.29697e-009, 1.30322e-009,
+ 1.30947e-009, 1.31572e-009, 1.32197e-009, 1.32822e-009)"
+          kdata_1to0_typ="(1, 0.969945, 0.967761, 0.965584, 0.963414, 0.961251,
+ 0.922663, 0.917876, 0.913122, 0.908402, 0.903714, 0.851047,
+ 0.843315, 0.835827, 0.828581, 0.821414, 0.777789, 0.768792,
+ 0.759918, 0.751166, 0.742532, 0.734016, 0.55307, 0.537138,
+ 0.52166, 0.506619, 0.491996, 0.366398, 0.350055, 0.334232,
+ 0.318906, 0.304052, 0.267484, 0.253148, 0.23932, 0.225815,
+ 0.212624, 0.239538, 0.228337, 0.217242, 0.206183, 0.204381,
+ 0.194033, 0.183877, 0.173777, 0.163736, 0.198952, 0.190664,
+ 0.182312, 0.1739, 0.165717, 0.170127, 0.16219, 0.154145,
+ 0.146131, 0.138011, 0.141711, 0.13341, 0.124857, 0.116071,
+ 0.107027, 0.153405, 0.145329, 0.136956, 0.128286, 0.11476,
+ 0.103503, 0.0919088, 0.0799865, 0.0670827, 0.0281211, 0.0117597,
+ 0, 0, 0, 0.0834382, 0.0701074, 0.0565091,
+ 0.0408893, 0.0245442, 0.0671925, 0.0543346, 0.0413051, 0.0277456,
+ 0.0127862, 0.00102775, 0, 0, 0, 0,
+ 0.0193647, 0.0104846, 0.00154843, 0, 0.0346995, 0.0293831,
+ 0.0239779, 0.0184849, 0.012905, 0.0133686, 0.00943205, 0.00530731,
+ 0.00108283, 0, 0.00937699, 0.00689617, 0.00437921, 0.00182603,
+ 0, 0.00216168, 0.000431909, 0, 0, 0,
+ 0.0182273, 0.0184874, 0.018742, 0.0189907, 0.0137603, 0.0140486,
+ 0.0143348, 0.014619, 0.0149012, 0.012462, 0.0127637, 0.0131749,
+ 0.0137195, 0.0142671, 0.00858316, 0.00888649, 0.00919061, 0.00949552,
+ 0.00980122, 0.00658873, 0.00668349, 0.00677755, 0.00687091, 0.00696356,
+ 0, 0, 0, 0, 0.0026533, 0.00305218,
+ 0.00345251, 0.00385433, 0.00425764, 0.00128215, 0.00147873, 0.0016757,
+ 0.00187306, 0.00207081, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0.00312929, 0.00354451, 0.00396081, 0.00437819, 0, 0,
+ 0, 0, 0, 0.00283054, 0.00324669, 0.00366393,
+ 0.00408225, 0.00450167, 0.00320158, 0.00351594, 0.00383091, 0.00414651,
+ 0.00446272, 0.00477956, 0.0034087, 0.00361956, 0.0038307, 0.00404212,
+ 0.00425382, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0.00147984,
+ 0.00168904, 0.00189851, 0.00210825, 0)"
+          vdata_typ="(-1.8, -1.74, -1.68, -1.62, -1.56, -1.5,
+ -1.44, -1.38, -1.32, -1.26, -1.2, -1.14,
+ -1.08, -1.02, -0.96, -0.9, -0.84, -0.78,
+ -0.72, -0.66, -0.6, -0.54, -0.48, -0.42,
+ -0.36, -0.3, -0.24, -0.18, -0.12, -0.06,
+ 0, 0.06, 0.12, 0.18, 0.24, 0.3,
+ 0.36, 0.42, 0.48, 0.54, 0.6, 0.66,
+ 0.72, 0.78, 0.84, 0.9, 0.96, 1.02,
+ 1.08, 1.14, 1.2, 1.26, 1.32, 1.38,
+ 1.44, 1.5, 1.56, 1.62, 1.68, 1.74,
+ 1.8, 1.86, 1.92, 1.98, 2.04, 2.1,
+ 2.16, 2.22, 2.28, 2.34, 2.4, 2.46,
+ 2.52, 2.58, 2.64, 2.7, 2.76, 2.82,
+ 2.88, 2.94, 3, 3.06, 3.12, 3.18,
+ 3.24, 3.3, 3.36, 3.42, 3.48, 3.54,
+ 3.6)"
+          idata_typ="(-6.345, -5.918, -5.492, -5.066, -4.64, -4.214,
+ -3.788, -3.363, -2.937, -2.511, -2.086, -1.663,
+ -1.243, -0.8341, -0.4448, -0.196, -0.1389, -0.1177,
+ -0.1018, -0.08764, -0.075, -0.06428, -0.05584, -0.04952,
+ -0.04448, -0.0399, -0.03541, -0.03094, -0.02644, -0.02194,
+ -0.01743, -0.01301, -0.008738, -0.004612, -0.0006315, 0.003204,
+ 0.006895, 0.01044, 0.01383, 0.01707, 0.02014, 0.02303,
+ 0.02573, 0.02821, 0.03045, 0.03244, 0.0342, 0.03576,
+ 0.03718, 0.03853, 0.03986, 0.0412, 0.04257, 0.04398,
+ 0.04543, 0.04695, 0.04854, 0.0502, 0.05195, 0.05377,
+ 0.05569, 0.0577, 0.05975, 0.06183, 0.06393, 0.06606,
+ 0.06826, 0.07067, 0.07359, 0.0773, 0.08184, 0.08709,
+ 0.09294, 0.09942, 0.1074, 0.1257, 0.2032, 0.3338,
+ 0.4821, 0.6392, 0.7982, 0.9575, 1.116, 1.276,
+ 1.435, 1.595, 1.754, 1.914, 2.073, 2.233,
+ 2.392)"
+          tdata_0to1_min="(1.63161e-011, 2.2246e-011, 2.81759e-011, 3.41058e-011, 4.00356e-011, 4.59655e-011,
+ 5.18954e-011, 5.78253e-011, 6.37551e-011, 6.9685e-011, 7.56149e-011, 8.15448e-011,
+ 8.74746e-011, 9.34045e-011, 9.93344e-011, 1.05264e-010, 1.11194e-010, 1.17124e-010,
+ 1.23054e-010, 1.28984e-010, 1.34914e-010, 1.40843e-010, 1.46773e-010, 1.52703e-010,
+ 1.58633e-010, 1.64563e-010, 1.70493e-010, 1.76423e-010, 1.82353e-010, 1.88282e-010,
+ 1.94212e-010, 2.00142e-010, 2.06072e-010, 2.12002e-010, 2.17932e-010, 2.23862e-010,
+ 2.29792e-010, 2.35721e-010, 2.41651e-010, 2.47581e-010, 2.53511e-010, 2.59441e-010,
+ 2.65371e-010, 2.71301e-010, 2.77231e-010, 2.8316e-010, 2.8909e-010, 2.9502e-010,
+ 3.0095e-010, 3.0688e-010, 3.1281e-010, 3.1874e-010, 3.2467e-010, 3.30599e-010,
+ 3.36529e-010, 3.42459e-010, 3.48389e-010, 3.54319e-010, 3.60249e-010, 3.66179e-010,
+ 3.72109e-010, 3.78038e-010, 3.83968e-010, 3.89898e-010, 3.95828e-010, 4.01758e-010,
+ 4.07688e-010, 4.13618e-010, 4.19548e-010, 4.25477e-010, 4.31407e-010, 4.37337e-010,
+ 4.43267e-010, 4.49197e-010, 4.55127e-010, 4.61057e-010, 4.66987e-010, 4.72916e-010,
+ 4.78846e-010, 4.84776e-010, 4.90706e-010, 4.96636e-010, 5.02566e-010, 5.08496e-010,
+ 5.14426e-010, 5.20355e-010, 5.26285e-010, 5.32215e-010, 5.38145e-010, 5.44075e-010,
+ 5.50005e-010, 5.55935e-010, 5.61865e-010, 5.67794e-010, 5.73724e-010, 5.79654e-010,
+ 5.85584e-010, 5.91514e-010, 5.97444e-010, 6.03374e-010, 6.09304e-010, 6.15233e-010,
+ 6.21163e-010, 6.27093e-010, 6.33023e-010, 6.38953e-010, 6.44883e-010, 6.50813e-010,
+ 6.56743e-010, 6.62672e-010, 6.68602e-010, 6.74532e-010, 6.80462e-010, 6.86392e-010,
+ 6.92322e-010, 6.98252e-010, 7.04182e-010, 7.10111e-010, 7.16041e-010, 7.21971e-010,
+ 7.27901e-010, 7.33831e-010, 7.39761e-010, 7.45691e-010, 7.51621e-010, 7.5755e-010,
+ 7.6348e-010, 7.6941e-010, 7.7534e-010, 7.8127e-010, 7.872e-010, 7.9313e-010,
+ 7.9906e-010, 8.04989e-010, 8.10919e-010, 8.16849e-010, 8.22779e-010, 8.28709e-010,
+ 8.34639e-010, 8.40569e-010, 8.46499e-010, 8.52428e-010, 8.58358e-010, 8.64288e-010,
+ 8.70218e-010, 8.76148e-010, 8.82078e-010, 8.88008e-010, 8.93938e-010, 8.99867e-010,
+ 9.05797e-010, 9.11727e-010, 9.17657e-010, 9.23587e-010, 9.29517e-010, 9.35447e-010,
+ 9.41377e-010, 9.47306e-010, 9.53236e-010, 9.59166e-010, 9.65096e-010, 9.71026e-010,
+ 9.76956e-010, 9.82886e-010, 9.88816e-010, 9.94745e-010, 1.00068e-009, 1.00661e-009,
+ 1.01254e-009, 1.01846e-009, 1.02439e-009, 1.03032e-009, 1.03625e-009, 1.04218e-009,
+ 1.04811e-009, 1.05404e-009, 1.05997e-009, 1.0659e-009, 1.07183e-009, 1.07776e-009,
+ 1.08369e-009, 1.08962e-009, 1.09555e-009, 1.10148e-009, 1.10741e-009, 1.11334e-009,
+ 1.11927e-009, 1.1252e-009, 1.13113e-009, 1.13706e-009, 1.14299e-009, 1.14892e-009,
+ 1.15485e-009, 1.16078e-009, 1.16671e-009, 1.17264e-009, 1.17857e-009, 1.1845e-009,
+ 1.19043e-009, 1.19636e-009, 1.20229e-009, 1.20822e-009)"
+          kdata_0to1_min="(0, 0.00693597, 0.00734267, 0.00775038, 0.00815913, 0.00858505,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0.0149774, 0.0168403, 0.0186985, 0.0205519,
+ 0.0224006, 0.0240851, 0.0257124, 0.0534193, 0.0575498, 0.0616171,
+ 0.0656214, 0.069563, 0.102944, 0.109289, 0.1155, 0.121575,
+ 0.127512, 0.185885, 0.194014, 0.201885, 0.209487, 0.216904,
+ 0.262763, 0.270595, 0.278029, 0.284935, 0.291331, 0.389536,
+ 0.397239, 0.403807, 0.409531, 0.41272, 0.458302, 0.460574,
+ 0.460332, 0.45866, 0.456168, 0.521521, 0.519402, 0.516554,
+ 0.512182, 0.507981, 0.562714, 0.560143, 0.557616, 0.556013,
+ 0.55331, 0.659015, 0.662791, 0.666581, 0.669294, 0.672524,
+ 0.716442, 0.724711, 0.731962, 0.740509, 0.749691, 0.739752,
+ 0.749267, 0.759439, 0.770012, 0.780565, 0.791097, 0.79587,
+ 0.809271, 0.822809, 0.836161, 0.849325, 0.834494, 0.847778,
+ 0.862015, 0.876457, 0.891109, 0.864523, 0.877546, 0.890758,
+ 0.904235, 0.918949, 0.917735, 0.932302, 0.946993, 0.961955,
+ 0.977195, 0.924242, 0.935102, 0.946108, 0.957264, 0.968572,
+ 0.909004, 0.915836, 0.922722, 0.929662, 0.936656, 0.952113,
+ 0.960445, 0.968871, 0.977393, 0.986011, 0.960073, 0.966314,
+ 0.972606, 0.97895, 0.985348, 0.970999, 0.976042, 0.98112,
+ 0.986232, 0.991379, 0.972387, 0.975803, 0.979234, 0.98268,
+ 0.986141, 0.967094, 0.968918, 0.970746, 0.972578, 0.974414,
+ 0.973267, 0.97489, 0.976515, 0.978144, 0.979776, 0.98008,
+ 0.981606, 0.983135, 0.984771, 0.986428, 0.984285, 0.985785,
+ 0.987287, 0.988793, 0.990302, 0.982654, 0.983469, 0.984284,
+ 0.9851, 0.985918, 0.989565, 0.990614, 0.991664, 0.992715,
+ 0.993768, 0.993327, 0.994265, 0.995205, 0.996146, 0.997089,
+ 0.998032, 1, 1, 1, 1, 1,
+ 0.99667, 0.997028, 0.997387, 0.997745, 0.998104, 0.993811,
+ 0.993821, 0.99383, 0.99384, 0.993849, 0.998489, 0.998848,
+ 0.999207, 0.999566, 0.999926, 0.998882, 0.999149, 0.999417,
+ 0.999684, 0.999951, 1, 1)"
+          tdata_1to0_min="(7.19709e-011, 7.82209e-011, 8.44709e-011, 9.07209e-011, 9.69709e-011, 1.03221e-010,
+ 1.09471e-010, 1.15721e-010, 1.21971e-010, 1.28221e-010, 1.34471e-010, 1.40721e-010,
+ 1.46971e-010, 1.53221e-010, 1.59471e-010, 1.65721e-010, 1.71971e-010, 1.78221e-010,
+ 1.84471e-010, 1.90721e-010, 1.96971e-010, 2.03221e-010, 2.09471e-010, 2.15721e-010,
+ 2.21971e-010, 2.28221e-010, 2.34471e-010, 2.40721e-010, 2.46971e-010, 2.53221e-010,
+ 2.59471e-010, 2.65721e-010, 2.71971e-010, 2.78221e-010, 2.84471e-010, 2.90721e-010,
+ 2.96971e-010, 3.03221e-010, 3.09471e-010, 3.15721e-010, 3.21971e-010, 3.28221e-010,
+ 3.34471e-010, 3.40721e-010, 3.46971e-010, 3.53221e-010, 3.59471e-010, 3.65721e-010,
+ 3.71971e-010, 3.78221e-010, 3.84471e-010, 3.90721e-010, 3.96971e-010, 4.03221e-010,
+ 4.09471e-010, 4.15721e-010, 4.21971e-010, 4.28221e-010, 4.34471e-010, 4.40721e-010,
+ 4.46971e-010, 4.53221e-010, 4.59471e-010, 4.65721e-010, 4.71971e-010, 4.78221e-010,
+ 4.84471e-010, 4.90721e-010, 4.96971e-010, 5.03221e-010, 5.09471e-010, 5.15721e-010,
+ 5.21971e-010, 5.28221e-010, 5.34471e-010, 5.40721e-010, 5.46971e-010, 5.53221e-010,
+ 5.59471e-010, 5.65721e-010, 5.71971e-010, 5.78221e-010, 5.84471e-010, 5.90721e-010,
+ 5.96971e-010, 6.03221e-010, 6.09471e-010, 6.15721e-010, 6.21971e-010, 6.28221e-010,
+ 6.34471e-010, 6.40721e-010, 6.46971e-010, 6.53221e-010, 6.59471e-010, 6.65721e-010,
+ 6.71971e-010, 6.78221e-010, 6.84471e-010, 6.90721e-010, 6.96971e-010, 7.03221e-010,
+ 7.09471e-010, 7.15721e-010, 7.21971e-010, 7.28221e-010, 7.34471e-010, 7.40721e-010,
+ 7.46971e-010, 7.53221e-010, 7.59471e-010, 7.65721e-010, 7.71971e-010, 7.78221e-010,
+ 7.84471e-010, 7.90721e-010, 7.96971e-010, 8.03221e-010, 8.09471e-010, 8.15721e-010,
+ 8.21971e-010, 8.28221e-010, 8.34471e-010, 8.40721e-010, 8.46971e-010, 8.53221e-010,
+ 8.59471e-010, 8.65721e-010, 8.71971e-010, 8.78221e-010, 8.84471e-010, 8.90721e-010,
+ 8.96971e-010, 9.03221e-010, 9.09471e-010, 9.15721e-010, 9.21971e-010, 9.28221e-010,
+ 9.34471e-010, 9.40721e-010, 9.46971e-010, 9.53221e-010, 9.59471e-010, 9.65721e-010,
+ 9.71971e-010, 9.78221e-010, 9.84471e-010, 9.90721e-010, 9.96971e-010, 1.00322e-009,
+ 1.00947e-009, 1.01572e-009, 1.02197e-009, 1.02822e-009, 1.03447e-009, 1.04072e-009,
+ 1.04697e-009, 1.05322e-009, 1.05947e-009, 1.06572e-009, 1.07197e-009, 1.07822e-009,
+ 1.08447e-009, 1.09072e-009, 1.09697e-009, 1.10322e-009, 1.10947e-009, 1.11572e-009,
+ 1.12197e-009, 1.12822e-009, 1.13447e-009, 1.14072e-009, 1.14697e-009, 1.15322e-009,
+ 1.15947e-009, 1.16572e-009, 1.17197e-009, 1.17822e-009, 1.18447e-009, 1.19072e-009,
+ 1.19697e-009, 1.20322e-009, 1.20947e-009, 1.21572e-009, 1.22197e-009, 1.22822e-009,
+ 1.23447e-009, 1.24072e-009, 1.24697e-009, 1.25322e-009, 1.25947e-009, 1.26572e-009,
+ 1.27197e-009, 1.27822e-009, 1.28447e-009, 1.29072e-009, 1.29697e-009, 1.30322e-009,
+ 1.30947e-009, 1.31572e-009, 1.32197e-009, 1.32822e-009)"
+          kdata_1to0_min="(1, 0.969945, 0.967761, 0.965584, 0.963414, 0.961251,
+ 0.922663, 0.917876, 0.913122, 0.908402, 0.903714, 0.851047,
+ 0.843315, 0.835827, 0.828581, 0.821414, 0.777789, 0.768792,
+ 0.759918, 0.751166, 0.742532, 0.734016, 0.55307, 0.537138,
+ 0.52166, 0.506619, 0.491996, 0.366398, 0.350055, 0.334232,
+ 0.318906, 0.304052, 0.267484, 0.253148, 0.23932, 0.225815,
+ 0.212624, 0.239538, 0.228337, 0.217242, 0.206183, 0.204381,
+ 0.194033, 0.183877, 0.173777, 0.163736, 0.198952, 0.190664,
+ 0.182312, 0.1739, 0.165717, 0.170127, 0.16219, 0.154145,
+ 0.146131, 0.138011, 0.141711, 0.13341, 0.124857, 0.116071,
+ 0.107027, 0.153405, 0.145329, 0.136956, 0.128286, 0.11476,
+ 0.103503, 0.0919088, 0.0799865, 0.0670827, 0.0281211, 0.0117597,
+ 0, 0, 0, 0.0834382, 0.0701074, 0.0565091,
+ 0.0408893, 0.0245442, 0.0671925, 0.0543346, 0.0413051, 0.0277456,
+ 0.0127862, 0.00102775, 0, 0, 0, 0,
+ 0.0193647, 0.0104846, 0.00154843, 0, 0.0346995, 0.0293831,
+ 0.0239779, 0.0184849, 0.012905, 0.0133686, 0.00943205, 0.00530731,
+ 0.00108283, 0, 0.00937699, 0.00689617, 0.00437921, 0.00182603,
+ 0, 0.00216168, 0.000431909, 0, 0, 0,
+ 0.0182273, 0.0184874, 0.018742, 0.0189907, 0.0137603, 0.0140486,
+ 0.0143348, 0.014619, 0.0149012, 0.012462, 0.0127637, 0.0131749,
+ 0.0137195, 0.0142671, 0.00858316, 0.00888649, 0.00919061, 0.00949552,
+ 0.00980122, 0.00658873, 0.00668349, 0.00677755, 0.00687091, 0.00696356,
+ 0, 0, 0, 0, 0.0026533, 0.00305218,
+ 0.00345251, 0.00385433, 0.00425764, 0.00128215, 0.00147873, 0.0016757,
+ 0.00187306, 0.00207081, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0.00312929, 0.00354451, 0.00396081, 0.00437819, 0, 0,
+ 0, 0, 0, 0.00283054, 0.00324669, 0.00366393,
+ 0.00408225, 0.00450167, 0.00320158, 0.00351594, 0.00383091, 0.00414651,
+ 0.00446272, 0.00477956, 0.0034087, 0.00361956, 0.0038307, 0.00404212,
+ 0.00425382, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0.00147984,
+ 0.00168904, 0.00189851, 0.00210825, 0)"
+          vdata_min="(-1.8, -1.74, -1.68, -1.62, -1.56, -1.5,
+ -1.44, -1.38, -1.32, -1.26, -1.2, -1.14,
+ -1.08, -1.02, -0.96, -0.9, -0.84, -0.78,
+ -0.72, -0.66, -0.6, -0.54, -0.48, -0.42,
+ -0.36, -0.3, -0.24, -0.18, -0.12, -0.06,
+ 0, 0.06, 0.12, 0.18, 0.24, 0.3,
+ 0.36, 0.42, 0.48, 0.54, 0.6, 0.66,
+ 0.72, 0.78, 0.84, 0.9, 0.96, 1.02,
+ 1.08, 1.14, 1.2, 1.26, 1.32, 1.38,
+ 1.44, 1.5, 1.56, 1.62, 1.68, 1.74,
+ 1.8, 1.86, 1.92, 1.98, 2.04, 2.1,
+ 2.16, 2.22, 2.28, 2.34, 2.4, 2.46,
+ 2.52, 2.58, 2.64, 2.7, 2.76, 2.82,
+ 2.88, 2.94, 3, 3.06, 3.12, 3.18,
+ 3.24, 3.3, 3.36, 3.42, 3.48, 3.54,
+ 3.6)"
+          idata_min="(-6.345, -5.918, -5.492, -5.066, -4.64, -4.214,
+ -3.788, -3.363, -2.937, -2.511, -2.086, -1.663,
+ -1.243, -0.8341, -0.4448, -0.196, -0.1389, -0.1177,
+ -0.1018, -0.08764, -0.075, -0.06428, -0.05584, -0.04952,
+ -0.04448, -0.0399, -0.03541, -0.03094, -0.02644, -0.02194,
+ -0.01743, -0.01301, -0.008738, -0.004612, -0.0006315, 0.003204,
+ 0.006895, 0.01044, 0.01383, 0.01707, 0.02014, 0.02303,
+ 0.02573, 0.02821, 0.03045, 0.03244, 0.0342, 0.03576,
+ 0.03718, 0.03853, 0.03986, 0.0412, 0.04257, 0.04398,
+ 0.04543, 0.04695, 0.04854, 0.0502, 0.05195, 0.05377,
+ 0.05569, 0.0577, 0.05975, 0.06183, 0.06393, 0.06606,
+ 0.06826, 0.07067, 0.07359, 0.0773, 0.08184, 0.08709,
+ 0.09294, 0.09942, 0.1074, 0.1257, 0.2032, 0.3338,
+ 0.4821, 0.6392, 0.7982, 0.9575, 1.116, 1.276,
+ 1.435, 1.595, 1.754, 1.914, 2.073, 2.233,
+ 2.392)"
+          tdata_0to1_max="(1.63161e-011, 2.2246e-011, 2.81759e-011, 3.41058e-011, 4.00356e-011, 4.59655e-011,
+ 5.18954e-011, 5.78253e-011, 6.37551e-011, 6.9685e-011, 7.56149e-011, 8.15448e-011,
+ 8.74746e-011, 9.34045e-011, 9.93344e-011, 1.05264e-010, 1.11194e-010, 1.17124e-010,
+ 1.23054e-010, 1.28984e-010, 1.34914e-010, 1.40843e-010, 1.46773e-010, 1.52703e-010,
+ 1.58633e-010, 1.64563e-010, 1.70493e-010, 1.76423e-010, 1.82353e-010, 1.88282e-010,
+ 1.94212e-010, 2.00142e-010, 2.06072e-010, 2.12002e-010, 2.17932e-010, 2.23862e-010,
+ 2.29792e-010, 2.35721e-010, 2.41651e-010, 2.47581e-010, 2.53511e-010, 2.59441e-010,
+ 2.65371e-010, 2.71301e-010, 2.77231e-010, 2.8316e-010, 2.8909e-010, 2.9502e-010,
+ 3.0095e-010, 3.0688e-010, 3.1281e-010, 3.1874e-010, 3.2467e-010, 3.30599e-010,
+ 3.36529e-010, 3.42459e-010, 3.48389e-010, 3.54319e-010, 3.60249e-010, 3.66179e-010,
+ 3.72109e-010, 3.78038e-010, 3.83968e-010, 3.89898e-010, 3.95828e-010, 4.01758e-010,
+ 4.07688e-010, 4.13618e-010, 4.19548e-010, 4.25477e-010, 4.31407e-010, 4.37337e-010,
+ 4.43267e-010, 4.49197e-010, 4.55127e-010, 4.61057e-010, 4.66987e-010, 4.72916e-010,
+ 4.78846e-010, 4.84776e-010, 4.90706e-010, 4.96636e-010, 5.02566e-010, 5.08496e-010,
+ 5.14426e-010, 5.20355e-010, 5.26285e-010, 5.32215e-010, 5.38145e-010, 5.44075e-010,
+ 5.50005e-010, 5.55935e-010, 5.61865e-010, 5.67794e-010, 5.73724e-010, 5.79654e-010,
+ 5.85584e-010, 5.91514e-010, 5.97444e-010, 6.03374e-010, 6.09304e-010, 6.15233e-010,
+ 6.21163e-010, 6.27093e-010, 6.33023e-010, 6.38953e-010, 6.44883e-010, 6.50813e-010,
+ 6.56743e-010, 6.62672e-010, 6.68602e-010, 6.74532e-010, 6.80462e-010, 6.86392e-010,
+ 6.92322e-010, 6.98252e-010, 7.04182e-010, 7.10111e-010, 7.16041e-010, 7.21971e-010,
+ 7.27901e-010, 7.33831e-010, 7.39761e-010, 7.45691e-010, 7.51621e-010, 7.5755e-010,
+ 7.6348e-010, 7.6941e-010, 7.7534e-010, 7.8127e-010, 7.872e-010, 7.9313e-010,
+ 7.9906e-010, 8.04989e-010, 8.10919e-010, 8.16849e-010, 8.22779e-010, 8.28709e-010,
+ 8.34639e-010, 8.40569e-010, 8.46499e-010, 8.52428e-010, 8.58358e-010, 8.64288e-010,
+ 8.70218e-010, 8.76148e-010, 8.82078e-010, 8.88008e-010, 8.93938e-010, 8.99867e-010,
+ 9.05797e-010, 9.11727e-010, 9.17657e-010, 9.23587e-010, 9.29517e-010, 9.35447e-010,
+ 9.41377e-010, 9.47306e-010, 9.53236e-010, 9.59166e-010, 9.65096e-010, 9.71026e-010,
+ 9.76956e-010, 9.82886e-010, 9.88816e-010, 9.94745e-010, 1.00068e-009, 1.00661e-009,
+ 1.01254e-009, 1.01846e-009, 1.02439e-009, 1.03032e-009, 1.03625e-009, 1.04218e-009,
+ 1.04811e-009, 1.05404e-009, 1.05997e-009, 1.0659e-009, 1.07183e-009, 1.07776e-009,
+ 1.08369e-009, 1.08962e-009, 1.09555e-009, 1.10148e-009, 1.10741e-009, 1.11334e-009,
+ 1.11927e-009, 1.1252e-009, 1.13113e-009, 1.13706e-009, 1.14299e-009, 1.14892e-009,
+ 1.15485e-009, 1.16078e-009, 1.16671e-009, 1.17264e-009, 1.17857e-009, 1.1845e-009,
+ 1.19043e-009, 1.19636e-009, 1.20229e-009, 1.20822e-009)"
+          kdata_0to1_max="(0, 0.00693597, 0.00734267, 0.00775038, 0.00815913, 0.00858505,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0.0149774, 0.0168403, 0.0186985, 0.0205519,
+ 0.0224006, 0.0240851, 0.0257124, 0.0534193, 0.0575498, 0.0616171,
+ 0.0656214, 0.069563, 0.102944, 0.109289, 0.1155, 0.121575,
+ 0.127512, 0.185885, 0.194014, 0.201885, 0.209487, 0.216904,
+ 0.262763, 0.270595, 0.278029, 0.284935, 0.291331, 0.389536,
+ 0.397239, 0.403807, 0.409531, 0.41272, 0.458302, 0.460574,
+ 0.460332, 0.45866, 0.456168, 0.521521, 0.519402, 0.516554,
+ 0.512182, 0.507981, 0.562714, 0.560143, 0.557616, 0.556013,
+ 0.55331, 0.659015, 0.662791, 0.666581, 0.669294, 0.672524,
+ 0.716442, 0.724711, 0.731962, 0.740509, 0.749691, 0.739752,
+ 0.749267, 0.759439, 0.770012, 0.780565, 0.791097, 0.79587,
+ 0.809271, 0.822809, 0.836161, 0.849325, 0.834494, 0.847778,
+ 0.862015, 0.876457, 0.891109, 0.864523, 0.877546, 0.890758,
+ 0.904235, 0.918949, 0.917735, 0.932302, 0.946993, 0.961955,
+ 0.977195, 0.924242, 0.935102, 0.946108, 0.957264, 0.968572,
+ 0.909004, 0.915836, 0.922722, 0.929662, 0.936656, 0.952113,
+ 0.960445, 0.968871, 0.977393, 0.986011, 0.960073, 0.966314,
+ 0.972606, 0.97895, 0.985348, 0.970999, 0.976042, 0.98112,
+ 0.986232, 0.991379, 0.972387, 0.975803, 0.979234, 0.98268,
+ 0.986141, 0.967094, 0.968918, 0.970746, 0.972578, 0.974414,
+ 0.973267, 0.97489, 0.976515, 0.978144, 0.979776, 0.98008,
+ 0.981606, 0.983135, 0.984771, 0.986428, 0.984285, 0.985785,
+ 0.987287, 0.988793, 0.990302, 0.982654, 0.983469, 0.984284,
+ 0.9851, 0.985918, 0.989565, 0.990614, 0.991664, 0.992715,
+ 0.993768, 0.993327, 0.994265, 0.995205, 0.996146, 0.997089,
+ 0.998032, 1, 1, 1, 1, 1,
+ 0.99667, 0.997028, 0.997387, 0.997745, 0.998104, 0.993811,
+ 0.993821, 0.99383, 0.99384, 0.993849, 0.998489, 0.998848,
+ 0.999207, 0.999566, 0.999926, 0.998882, 0.999149, 0.999417,
+ 0.999684, 0.999951, 1, 1)"
+          tdata_1to0_max="(7.19709e-011, 7.82209e-011, 8.44709e-011, 9.07209e-011, 9.69709e-011, 1.03221e-010,
+ 1.09471e-010, 1.15721e-010, 1.21971e-010, 1.28221e-010, 1.34471e-010, 1.40721e-010,
+ 1.46971e-010, 1.53221e-010, 1.59471e-010, 1.65721e-010, 1.71971e-010, 1.78221e-010,
+ 1.84471e-010, 1.90721e-010, 1.96971e-010, 2.03221e-010, 2.09471e-010, 2.15721e-010,
+ 2.21971e-010, 2.28221e-010, 2.34471e-010, 2.40721e-010, 2.46971e-010, 2.53221e-010,
+ 2.59471e-010, 2.65721e-010, 2.71971e-010, 2.78221e-010, 2.84471e-010, 2.90721e-010,
+ 2.96971e-010, 3.03221e-010, 3.09471e-010, 3.15721e-010, 3.21971e-010, 3.28221e-010,
+ 3.34471e-010, 3.40721e-010, 3.46971e-010, 3.53221e-010, 3.59471e-010, 3.65721e-010,
+ 3.71971e-010, 3.78221e-010, 3.84471e-010, 3.90721e-010, 3.96971e-010, 4.03221e-010,
+ 4.09471e-010, 4.15721e-010, 4.21971e-010, 4.28221e-010, 4.34471e-010, 4.40721e-010,
+ 4.46971e-010, 4.53221e-010, 4.59471e-010, 4.65721e-010, 4.71971e-010, 4.78221e-010,
+ 4.84471e-010, 4.90721e-010, 4.96971e-010, 5.03221e-010, 5.09471e-010, 5.15721e-010,
+ 5.21971e-010, 5.28221e-010, 5.34471e-010, 5.40721e-010, 5.46971e-010, 5.53221e-010,
+ 5.59471e-010, 5.65721e-010, 5.71971e-010, 5.78221e-010, 5.84471e-010, 5.90721e-010,
+ 5.96971e-010, 6.03221e-010, 6.09471e-010, 6.15721e-010, 6.21971e-010, 6.28221e-010,
+ 6.34471e-010, 6.40721e-010, 6.46971e-010, 6.53221e-010, 6.59471e-010, 6.65721e-010,
+ 6.71971e-010, 6.78221e-010, 6.84471e-010, 6.90721e-010, 6.96971e-010, 7.03221e-010,
+ 7.09471e-010, 7.15721e-010, 7.21971e-010, 7.28221e-010, 7.34471e-010, 7.40721e-010,
+ 7.46971e-010, 7.53221e-010, 7.59471e-010, 7.65721e-010, 7.71971e-010, 7.78221e-010,
+ 7.84471e-010, 7.90721e-010, 7.96971e-010, 8.03221e-010, 8.09471e-010, 8.15721e-010,
+ 8.21971e-010, 8.28221e-010, 8.34471e-010, 8.40721e-010, 8.46971e-010, 8.53221e-010,
+ 8.59471e-010, 8.65721e-010, 8.71971e-010, 8.78221e-010, 8.84471e-010, 8.90721e-010,
+ 8.96971e-010, 9.03221e-010, 9.09471e-010, 9.15721e-010, 9.21971e-010, 9.28221e-010,
+ 9.34471e-010, 9.40721e-010, 9.46971e-010, 9.53221e-010, 9.59471e-010, 9.65721e-010,
+ 9.71971e-010, 9.78221e-010, 9.84471e-010, 9.90721e-010, 9.96971e-010, 1.00322e-009,
+ 1.00947e-009, 1.01572e-009, 1.02197e-009, 1.02822e-009, 1.03447e-009, 1.04072e-009,
+ 1.04697e-009, 1.05322e-009, 1.05947e-009, 1.06572e-009, 1.07197e-009, 1.07822e-009,
+ 1.08447e-009, 1.09072e-009, 1.09697e-009, 1.10322e-009, 1.10947e-009, 1.11572e-009,
+ 1.12197e-009, 1.12822e-009, 1.13447e-009, 1.14072e-009, 1.14697e-009, 1.15322e-009,
+ 1.15947e-009, 1.16572e-009, 1.17197e-009, 1.17822e-009, 1.18447e-009, 1.19072e-009,
+ 1.19697e-009, 1.20322e-009, 1.20947e-009, 1.21572e-009, 1.22197e-009, 1.22822e-009,
+ 1.23447e-009, 1.24072e-009, 1.24697e-009, 1.25322e-009, 1.25947e-009, 1.26572e-009,
+ 1.27197e-009, 1.27822e-009, 1.28447e-009, 1.29072e-009, 1.29697e-009, 1.30322e-009,
+ 1.30947e-009, 1.31572e-009, 1.32197e-009, 1.32822e-009)"
+          kdata_1to0_max="(1, 0.969945, 0.967761, 0.965584, 0.963414, 0.961251,
+ 0.922663, 0.917876, 0.913122, 0.908402, 0.903714, 0.851047,
+ 0.843315, 0.835827, 0.828581, 0.821414, 0.777789, 0.768792,
+ 0.759918, 0.751166, 0.742532, 0.734016, 0.55307, 0.537138,
+ 0.52166, 0.506619, 0.491996, 0.366398, 0.350055, 0.334232,
+ 0.318906, 0.304052, 0.267484, 0.253148, 0.23932, 0.225815,
+ 0.212624, 0.239538, 0.228337, 0.217242, 0.206183, 0.204381,
+ 0.194033, 0.183877, 0.173777, 0.163736, 0.198952, 0.190664,
+ 0.182312, 0.1739, 0.165717, 0.170127, 0.16219, 0.154145,
+ 0.146131, 0.138011, 0.141711, 0.13341, 0.124857, 0.116071,
+ 0.107027, 0.153405, 0.145329, 0.136956, 0.128286, 0.11476,
+ 0.103503, 0.0919088, 0.0799865, 0.0670827, 0.0281211, 0.0117597,
+ 0, 0, 0, 0.0834382, 0.0701074, 0.0565091,
+ 0.0408893, 0.0245442, 0.0671925, 0.0543346, 0.0413051, 0.0277456,
+ 0.0127862, 0.00102775, 0, 0, 0, 0,
+ 0.0193647, 0.0104846, 0.00154843, 0, 0.0346995, 0.0293831,
+ 0.0239779, 0.0184849, 0.012905, 0.0133686, 0.00943205, 0.00530731,
+ 0.00108283, 0, 0.00937699, 0.00689617, 0.00437921, 0.00182603,
+ 0, 0.00216168, 0.000431909, 0, 0, 0,
+ 0.0182273, 0.0184874, 0.018742, 0.0189907, 0.0137603, 0.0140486,
+ 0.0143348, 0.014619, 0.0149012, 0.012462, 0.0127637, 0.0131749,
+ 0.0137195, 0.0142671, 0.00858316, 0.00888649, 0.00919061, 0.00949552,
+ 0.00980122, 0.00658873, 0.00668349, 0.00677755, 0.00687091, 0.00696356,
+ 0, 0, 0, 0, 0.0026533, 0.00305218,
+ 0.00345251, 0.00385433, 0.00425764, 0.00128215, 0.00147873, 0.0016757,
+ 0.00187306, 0.00207081, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0.00312929, 0.00354451, 0.00396081, 0.00437819, 0, 0,
+ 0, 0, 0, 0.00283054, 0.00324669, 0.00366393,
+ 0.00408225, 0.00450167, 0.00320158, 0.00351594, 0.00383091, 0.00414651,
+ 0.00446272, 0.00477956, 0.0034087, 0.00361956, 0.0038307, 0.00404212,
+ 0.00425382, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0.00147984,
+ 0.00168904, 0.00189851, 0.00210825, 0)"
+          vdata_max="(-1.8, -1.74, -1.68, -1.62, -1.56, -1.5,
+ -1.44, -1.38, -1.32, -1.26, -1.2, -1.14,
+ -1.08, -1.02, -0.96, -0.9, -0.84, -0.78,
+ -0.72, -0.66, -0.6, -0.54, -0.48, -0.42,
+ -0.36, -0.3, -0.24, -0.18, -0.12, -0.06,
+ 0, 0.06, 0.12, 0.18, 0.24, 0.3,
+ 0.36, 0.42, 0.48, 0.54, 0.6, 0.66,
+ 0.72, 0.78, 0.84, 0.9, 0.96, 1.02,
+ 1.08, 1.14, 1.2, 1.26, 1.32, 1.38,
+ 1.44, 1.5, 1.56, 1.62, 1.68, 1.74,
+ 1.8, 1.86, 1.92, 1.98, 2.04, 2.1,
+ 2.16, 2.22, 2.28, 2.34, 2.4, 2.46,
+ 2.52, 2.58, 2.64, 2.7, 2.76, 2.82,
+ 2.88, 2.94, 3, 3.06, 3.12, 3.18,
+ 3.24, 3.3, 3.36, 3.42, 3.48, 3.54,
+ 3.6)"
+          idata_max="(-6.345, -5.918, -5.492, -5.066, -4.64, -4.214,
+ -3.788, -3.363, -2.937, -2.511, -2.086, -1.663,
+ -1.243, -0.8341, -0.4448, -0.196, -0.1389, -0.1177,
+ -0.1018, -0.08764, -0.075, -0.06428, -0.05584, -0.04952,
+ -0.04448, -0.0399, -0.03541, -0.03094, -0.02644, -0.02194,
+ -0.01743, -0.01301, -0.008738, -0.004612, -0.0006315, 0.003204,
+ 0.006895, 0.01044, 0.01383, 0.01707, 0.02014, 0.02303,
+ 0.02573, 0.02821, 0.03045, 0.03244, 0.0342, 0.03576,
+ 0.03718, 0.03853, 0.03986, 0.0412, 0.04257, 0.04398,
+ 0.04543, 0.04695, 0.04854, 0.0502, 0.05195, 0.05377,
+ 0.05569, 0.0577, 0.05975, 0.06183, 0.06393, 0.06606,
+ 0.06826, 0.07067, 0.07359, 0.0773, 0.08184, 0.08709,
+ 0.09294, 0.09942, 0.1074, 0.1257, 0.2032, 0.3338,
+ 0.4821, 0.6392, 0.7982, 0.9575, 1.116, 1.276,
+ 1.435, 1.595, 1.754, 1.914, 2.073, 2.233,
+ 2.392)"
+ PORT: a_PdRef
+       a_signal
+       d_pulldown_control


*IBIS Pullup tables
Y_PullUp ibis_ktiv(icx_behavioral)
+ GENERIC: corner="ibis_typ"
+          tdata_0to1_typ="(7.19709e-011, 7.82209e-011, 8.44709e-011, 9.07209e-011, 9.69709e-011, 1.03221e-010,
+ 1.09471e-010, 1.15721e-010, 1.21971e-010, 1.28221e-010, 1.34471e-010, 1.40721e-010,
+ 1.46971e-010, 1.53221e-010, 1.59471e-010, 1.65721e-010, 1.71971e-010, 1.78221e-010,
+ 1.84471e-010, 1.90721e-010, 1.96971e-010, 2.03221e-010, 2.09471e-010, 2.15721e-010,
+ 2.21971e-010, 2.28221e-010, 2.34471e-010, 2.40721e-010, 2.46971e-010, 2.53221e-010,
+ 2.59471e-010, 2.65721e-010, 2.71971e-010, 2.78221e-010, 2.84471e-010, 2.90721e-010,
+ 2.96971e-010, 3.03221e-010, 3.09471e-010, 3.15721e-010, 3.21971e-010, 3.28221e-010,
+ 3.34471e-010, 3.40721e-010, 3.46971e-010, 3.53221e-010, 3.59471e-010, 3.65721e-010,
+ 3.71971e-010, 3.78221e-010, 3.84471e-010, 3.90721e-010, 3.96971e-010, 4.03221e-010,
+ 4.09471e-010, 4.15721e-010, 4.21971e-010, 4.28221e-010, 4.34471e-010, 4.40721e-010,
+ 4.46971e-010, 4.53221e-010, 4.59471e-010, 4.65721e-010, 4.71971e-010, 4.78221e-010,
+ 4.84471e-010, 4.90721e-010, 4.96971e-010, 5.03221e-010, 5.09471e-010, 5.15721e-010,
+ 5.21971e-010, 5.28221e-010, 5.34471e-010, 5.40721e-010, 5.46971e-010, 5.53221e-010,
+ 5.59471e-010, 5.65721e-010, 5.71971e-010, 5.78221e-010, 5.84471e-010, 5.90721e-010,
+ 5.96971e-010, 6.03221e-010, 6.09471e-010, 6.15721e-010, 6.21971e-010, 6.28221e-010,
+ 6.34471e-010, 6.40721e-010, 6.46971e-010, 6.53221e-010, 6.59471e-010, 6.65721e-010,
+ 6.71971e-010, 6.78221e-010, 6.84471e-010, 6.90721e-010, 6.96971e-010, 7.03221e-010,
+ 7.09471e-010, 7.15721e-010, 7.21971e-010, 7.28221e-010, 7.34471e-010, 7.40721e-010,
+ 7.46971e-010, 7.53221e-010, 7.59471e-010, 7.65721e-010, 7.71971e-010, 7.78221e-010,
+ 7.84471e-010, 7.90721e-010, 7.96971e-010, 8.03221e-010, 8.09471e-010, 8.15721e-010,
+ 8.21971e-010, 8.28221e-010, 8.34471e-010, 8.40721e-010, 8.46971e-010, 8.53221e-010,
+ 8.59471e-010, 8.65721e-010, 8.71971e-010, 8.78221e-010, 8.84471e-010, 8.90721e-010,
+ 8.96971e-010, 9.03221e-010, 9.09471e-010, 9.15721e-010, 9.21971e-010, 9.28221e-010,
+ 9.34471e-010, 9.40721e-010, 9.46971e-010, 9.53221e-010, 9.59471e-010, 9.65721e-010,
+ 9.71971e-010, 9.78221e-010, 9.84471e-010, 9.90721e-010, 9.96971e-010, 1.00322e-009,
+ 1.00947e-009, 1.01572e-009, 1.02197e-009, 1.02822e-009, 1.03447e-009, 1.04072e-009,
+ 1.04697e-009, 1.05322e-009, 1.05947e-009, 1.06572e-009, 1.07197e-009, 1.07822e-009,
+ 1.08447e-009, 1.09072e-009, 1.09697e-009, 1.10322e-009, 1.10947e-009, 1.11572e-009,
+ 1.12197e-009, 1.12822e-009, 1.13447e-009, 1.14072e-009, 1.14697e-009, 1.15322e-009,
+ 1.15947e-009, 1.16572e-009, 1.17197e-009, 1.17822e-009, 1.18447e-009, 1.19072e-009,
+ 1.19697e-009, 1.20322e-009, 1.20947e-009, 1.21572e-009, 1.22197e-009, 1.22822e-009,
+ 1.23447e-009, 1.24072e-009, 1.24697e-009, 1.25322e-009, 1.25947e-009, 1.26572e-009,
+ 1.27197e-009, 1.27822e-009, 1.28447e-009, 1.29072e-009, 1.29697e-009, 1.30322e-009,
+ 1.30947e-009, 1.31572e-009, 1.32197e-009, 1.32822e-009)"
+          kdata_0to1_typ="(0, 0.00144844, 0.00161591, 0.00178283, 0.00194921, 0.00211506,
+ 0.0087038, 0.00937234, 0.0100361, 0.0106951, 0.0113493, 0.0221732,
+ 0.0235462, 0.0248913, 0.0262091, 0.027512, 0.0384896, 0.040387,
+ 0.0422566, 0.0440992, 0.0459152, 0.0477052, 0.0909226, 0.0947716,
+ 0.0985008, 0.102115, 0.10562, 0.151672, 0.156561, 0.161263,
+ 0.165788, 0.170143, 0.231451, 0.237879, 0.244041, 0.249991,
+ 0.255738, 0.306646, 0.314487, 0.322133, 0.329544, 0.346723,
+ 0.354268, 0.361647, 0.368849, 0.375871, 0.436727, 0.446473,
+ 0.456075, 0.465528, 0.47489, 0.508024, 0.518296, 0.528421,
+ 0.538431, 0.548284, 0.578952, 0.589365, 0.599555, 0.609511,
+ 0.619187, 0.661993, 0.673295, 0.684356, 0.695153, 0.695174,
+ 0.703634, 0.711667, 0.719248, 0.725866, 0.705895, 0.708557,
+ 0.710598, 0.711564, 0.710588, 0.813801, 0.819259, 0.824199,
+ 0.827163, 0.82912, 0.854347, 0.858385, 0.861996, 0.865003,
+ 0.86646, 0.82184, 0.821897, 0.821674, 0.821592, 0.821429,
+ 0.86842, 0.871631, 0.874676, 0.877554, 0.928498, 0.936229,
+ 0.943903, 0.951517, 0.95907, 0.902802, 0.908617, 0.914903,
+ 0.921194, 0.927466, 0.912617, 0.919099, 0.925592, 0.932094,
+ 0.938605, 0.915914, 0.921739, 0.928803, 0.935927, 0.943095,
+ 0.982139, 0.992066, 1, 1, 0.970056, 0.977633,
+ 0.985279, 0.992996, 1, 0.981505, 0.988024, 0.995008,
+ 1, 1, 0.97652, 0.981778, 0.987072, 0.992403,
+ 0.997772, 0.989569, 0.994141, 0.99874, 1, 1,
+ 0.958503, 0.959695, 0.960888, 0.961952, 0.984313, 0.987439,
+ 0.99058, 0.993734, 0.996902, 0.986424, 0.988754, 0.991091,
+ 0.993435, 0.995786, 0.984205, 0.985709, 0.987216, 0.988726,
+ 0.990238, 0.991754, 0.993272, 0.994792, 0.996316, 0.997843,
+ 0.997771, 0.99948, 1, 1, 0.978729, 0.978557,
+ 0.978385, 0.978213, 0.978042, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 0.984196, 0.983159, 0.982125, 0.981093, 0.980062,
+ 0.991678, 0.991678, 0.991678, 0.991678, 0.991678, 1,
+ 1, 1, 1, 1)"
+          tdata_1to0_typ="(1.63161e-011, 2.2246e-011, 2.81759e-011, 3.41058e-011, 4.00356e-011, 4.59655e-011,
+ 5.18954e-011, 5.78253e-011, 6.37551e-011, 6.9685e-011, 7.56149e-011, 8.15448e-011,
+ 8.74746e-011, 9.34045e-011, 9.93344e-011, 1.05264e-010, 1.11194e-010, 1.17124e-010,
+ 1.23054e-010, 1.28984e-010, 1.34914e-010, 1.40843e-010, 1.46773e-010, 1.52703e-010,
+ 1.58633e-010, 1.64563e-010, 1.70493e-010, 1.76423e-010, 1.82353e-010, 1.88282e-010,
+ 1.94212e-010, 2.00142e-010, 2.06072e-010, 2.12002e-010, 2.17932e-010, 2.23862e-010,
+ 2.29792e-010, 2.35721e-010, 2.41651e-010, 2.47581e-010, 2.53511e-010, 2.59441e-010,
+ 2.65371e-010, 2.71301e-010, 2.77231e-010, 2.8316e-010, 2.8909e-010, 2.9502e-010,
+ 3.0095e-010, 3.0688e-010, 3.1281e-010, 3.1874e-010, 3.2467e-010, 3.30599e-010,
+ 3.36529e-010, 3.42459e-010, 3.48389e-010, 3.54319e-010, 3.60249e-010, 3.66179e-010,
+ 3.72109e-010, 3.78038e-010, 3.83968e-010, 3.89898e-010, 3.95828e-010, 4.01758e-010,
+ 4.07688e-010, 4.13618e-010, 4.19548e-010, 4.25477e-010, 4.31407e-010, 4.37337e-010,
+ 4.43267e-010, 4.49197e-010, 4.55127e-010, 4.61057e-010, 4.66987e-010, 4.72916e-010,
+ 4.78846e-010, 4.84776e-010, 4.90706e-010, 4.96636e-010, 5.02566e-010, 5.08496e-010,
+ 5.14426e-010, 5.20355e-010, 5.26285e-010, 5.32215e-010, 5.38145e-010, 5.44075e-010,
+ 5.50005e-010, 5.55935e-010, 5.61865e-010, 5.67794e-010, 5.73724e-010, 5.79654e-010,
+ 5.85584e-010, 5.91514e-010, 5.97444e-010, 6.03374e-010, 6.09304e-010, 6.15233e-010,
+ 6.21163e-010, 6.27093e-010, 6.33023e-010, 6.38953e-010, 6.44883e-010, 6.50813e-010,
+ 6.56743e-010, 6.62672e-010, 6.68602e-010, 6.74532e-010, 6.80462e-010, 6.86392e-010,
+ 6.92322e-010, 6.98252e-010, 7.04182e-010, 7.10111e-010, 7.16041e-010, 7.21971e-010,
+ 7.27901e-010, 7.33831e-010, 7.39761e-010, 7.45691e-010, 7.51621e-010, 7.5755e-010,
+ 7.6348e-010, 7.6941e-010, 7.7534e-010, 7.8127e-010, 7.872e-010, 7.9313e-010,
+ 7.9906e-010, 8.04989e-010, 8.10919e-010, 8.16849e-010, 8.22779e-010, 8.28709e-010,
+ 8.34639e-010, 8.40569e-010, 8.46499e-010, 8.52428e-010, 8.58358e-010, 8.64288e-010,
+ 8.70218e-010, 8.76148e-010, 8.82078e-010, 8.88008e-010, 8.93938e-010, 8.99867e-010,
+ 9.05797e-010, 9.11727e-010, 9.17657e-010, 9.23587e-010, 9.29517e-010, 9.35447e-010,
+ 9.41377e-010, 9.47306e-010, 9.53236e-010, 9.59166e-010, 9.65096e-010, 9.71026e-010,
+ 9.76956e-010, 9.82886e-010, 9.88816e-010, 9.94745e-010, 1.00068e-009, 1.00661e-009,
+ 1.01254e-009, 1.01846e-009, 1.02439e-009, 1.03032e-009, 1.03625e-009, 1.04218e-009,
+ 1.04811e-009, 1.05404e-009, 1.05997e-009, 1.0659e-009, 1.07183e-009, 1.07776e-009,
+ 1.08369e-009, 1.08962e-009, 1.09555e-009, 1.10148e-009, 1.10741e-009, 1.11334e-009,
+ 1.11927e-009, 1.1252e-009, 1.13113e-009, 1.13706e-009, 1.14299e-009, 1.14892e-009,
+ 1.15485e-009, 1.16078e-009, 1.16671e-009, 1.17264e-009, 1.17857e-009, 1.1845e-009,
+ 1.19043e-009, 1.19636e-009, 1.20229e-009, 1.20822e-009)"
+          kdata_1to0_typ="(1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 0.944958, 0.941817, 0.939014,
+ 0.936329, 0.933652, 0.928097, 0.926197, 0.924296, 0.922394,
+ 0.920489, 0.918327, 0.916081, 0.742328, 0.734287, 0.726279,
+ 0.718306, 0.710366, 0.5818, 0.572814, 0.563786, 0.554718,
+ 0.545614, 0.432759, 0.422287, 0.411632, 0.400804, 0.390031,
+ 0.357675, 0.345405, 0.33285, 0.319786, 0.306318, 0.299028,
+ 0.281999, 0.263834, 0.245179, 0.224, 0.21373, 0.19043,
+ 0.164822, 0.138767, 0.11283, 0.168453, 0.142421, 0.11653,
+ 0.0898447, 0.064093, 0.12499, 0.101151, 0.0779349, 0.0556811,
+ 0.0329568, 0.116942, 0.0977118, 0.0785584, 0.0587776, 0.0393621,
+ 0.100619, 0.0856291, 0.0698708, 0.0543328, 0.0388455, 0.0738995,
+ 0.0617298, 0.0492707, 0.0366203, 0.0238299, 0.0109021, 0.0561065,
+ 0.0467763, 0.0372812, 0.0274446, 0.0172799, 0.0457196, 0.0381295,
+ 0.0304268, 0.0225745, 0.0145697, 0.0383468, 0.0325389, 0.0266255,
+ 0.0206042, 0.0144643, 0.0365308, 0.0322321, 0.0277894, 0.0232542,
+ 0.0186239, 0.028672, 0.025203, 0.0216809, 0.0181047, 0.0144733,
+ 0.0148853, 0.0116153, 0.00831567, 0.00498609, 0.0016262, 0.0188761,
+ 0.0170186, 0.015139, 0.0132368, 0.0113117, 0.0155086, 0.0140556,
+ 0.0125899, 0.0111111, 0.00961925, 0.0139533, 0.0129102, 0.0118597,
+ 0.0108016, 0.00973602, 0.0114324, 0.0105801, 0.00972376, 0.00886338,
+ 0.00799891, 0.00901914, 0.00830074, 0.00758063, 0.0068588, 0.00613525,
+ 0.00561266, 0.00490209, 0.00419006, 0.00347656, 0.00276158, 0.00173159,
+ 0.000988725, 0.000244458, 0, 0, 0.00391781, 0.00364127,
+ 0.00336415, 0.00308644, 0.00280814, 0.00360153, 0.003408, 0.00321424,
+ 0.00302027, 0.00282607, 0.00282379, 0.00264561, 0.00246717, 0.00228846,
+ 0.00210949, 0.00204093, 0.00187022, 0.00169929, 0.00152814, 0.00135675,
+ 0.00118514, 0.00121595, 0.00106019, 0.000904174, 0.000747895, 0.000591352,
+ 0.00127719, 0.00118284, 0.00108844, 0.000993996, 0.000899505, 0.000727513,
+ 0.000625664, 0.000523821, 0.000421982, 0.000320148, 0.000293503, 0.000198808,
+ 0.000104067, 9.27975e-006, 0, 0.0004531, 0.000407536, 0.000361956,
+ 0.000316359, 0.000270744, 0.000225112, 0)"
+          vdata_typ="(-1.8, -1.74, -1.68, -1.62, -1.56, -1.5,
+ -1.44, -1.38, -1.32, -1.26, -1.2, -1.14,
+ -1.08, -1.02, -0.96, -0.9, -0.84, -0.78,
+ -0.72, -0.66, -0.6, -0.54, -0.48, -0.42,
+ -0.36, -0.3, -0.24, -0.18, -0.12, -0.06,
+ 0, 0.06, 0.12, 0.18, 0.24, 0.3,
+ 0.36, 0.42, 0.48, 0.54, 0.6, 0.66,
+ 0.72, 0.78, 0.84, 0.9, 0.96, 1.02,
+ 1.08, 1.14, 1.2, 1.26, 1.32, 1.38,
+ 1.44, 1.5, 1.56, 1.62, 1.68, 1.74,
+ 1.8, 1.86, 1.92, 1.98, 2.04, 2.1,
+ 2.16, 2.22, 2.28, 2.34, 2.4, 2.46,
+ 2.52, 2.58, 2.64, 2.7, 2.76, 2.82,
+ 2.88, 2.94, 3, 3.06, 3.12, 3.18,
+ 3.24, 3.3, 3.36, 3.42, 3.48, 3.54,
+ 3.6)"
+          idata_typ="(-2.394, -2.235, -2.075, -1.915, -1.756, -1.596,
+ -1.437, -1.277, -1.118, -0.9586, -0.7993, -0.6403,
+ -0.4841, -0.3375, -0.2096, -0.1333, -0.1135, -0.1032,
+ -0.09427, -0.08574, -0.07761, -0.06996, -0.06286, -0.05631,
+ -0.05017, -0.04422, -0.03837, -0.03258, -0.02687, -0.02127,
+ -0.01578, -0.01053, -0.005574, -0.0009032, 0.003482, 0.007583,
+ 0.0114, 0.01494, 0.0182, 0.02119, 0.0239, 0.02632,
+ 0.02844, 0.03027, 0.03189, 0.03338, 0.03481, 0.0362,
+ 0.03759, 0.03898, 0.04039, 0.04181, 0.04324, 0.0447,
+ 0.04617, 0.04766, 0.04918, 0.05073, 0.0523, 0.0539,
+ 0.05554, 0.05721, 0.05887, 0.06051, 0.06215, 0.06379,
+ 0.06553, 0.06774, 0.07132, 0.07727, 0.08581, 0.09653,
+ 0.109, 0.1233, 0.143, 0.1988, 0.4466, 0.8356,
+ 1.244, 1.664, 2.088, 2.513, 2.938, 3.364,
+ 3.79, 4.216, 4.641, 5.067, 5.493, 5.919,
+ 6.346)"
+          tdata_0to1_min="(7.19709e-011, 7.82209e-011, 8.44709e-011, 9.07209e-011, 9.69709e-011, 1.03221e-010,
+ 1.09471e-010, 1.15721e-010, 1.21971e-010, 1.28221e-010, 1.34471e-010, 1.40721e-010,
+ 1.46971e-010, 1.53221e-010, 1.59471e-010, 1.65721e-010, 1.71971e-010, 1.78221e-010,
+ 1.84471e-010, 1.90721e-010, 1.96971e-010, 2.03221e-010, 2.09471e-010, 2.15721e-010,
+ 2.21971e-010, 2.28221e-010, 2.34471e-010, 2.40721e-010, 2.46971e-010, 2.53221e-010,
+ 2.59471e-010, 2.65721e-010, 2.71971e-010, 2.78221e-010, 2.84471e-010, 2.90721e-010,
+ 2.96971e-010, 3.03221e-010, 3.09471e-010, 3.15721e-010, 3.21971e-010, 3.28221e-010,
+ 3.34471e-010, 3.40721e-010, 3.46971e-010, 3.53221e-010, 3.59471e-010, 3.65721e-010,
+ 3.71971e-010, 3.78221e-010, 3.84471e-010, 3.90721e-010, 3.96971e-010, 4.03221e-010,
+ 4.09471e-010, 4.15721e-010, 4.21971e-010, 4.28221e-010, 4.34471e-010, 4.40721e-010,
+ 4.46971e-010, 4.53221e-010, 4.59471e-010, 4.65721e-010, 4.71971e-010, 4.78221e-010,
+ 4.84471e-010, 4.90721e-010, 4.96971e-010, 5.03221e-010, 5.09471e-010, 5.15721e-010,
+ 5.21971e-010, 5.28221e-010, 5.34471e-010, 5.40721e-010, 5.46971e-010, 5.53221e-010,
+ 5.59471e-010, 5.65721e-010, 5.71971e-010, 5.78221e-010, 5.84471e-010, 5.90721e-010,
+ 5.96971e-010, 6.03221e-010, 6.09471e-010, 6.15721e-010, 6.21971e-010, 6.28221e-010,
+ 6.34471e-010, 6.40721e-010, 6.46971e-010, 6.53221e-010, 6.59471e-010, 6.65721e-010,
+ 6.71971e-010, 6.78221e-010, 6.84471e-010, 6.90721e-010, 6.96971e-010, 7.03221e-010,
+ 7.09471e-010, 7.15721e-010, 7.21971e-010, 7.28221e-010, 7.34471e-010, 7.40721e-010,
+ 7.46971e-010, 7.53221e-010, 7.59471e-010, 7.65721e-010, 7.71971e-010, 7.78221e-010,
+ 7.84471e-010, 7.90721e-010, 7.96971e-010, 8.03221e-010, 8.09471e-010, 8.15721e-010,
+ 8.21971e-010, 8.28221e-010, 8.34471e-010, 8.40721e-010, 8.46971e-010, 8.53221e-010,
+ 8.59471e-010, 8.65721e-010, 8.71971e-010, 8.78221e-010, 8.84471e-010, 8.90721e-010,
+ 8.96971e-010, 9.03221e-010, 9.09471e-010, 9.15721e-010, 9.21971e-010, 9.28221e-010,
+ 9.34471e-010, 9.40721e-010, 9.46971e-010, 9.53221e-010, 9.59471e-010, 9.65721e-010,
+ 9.71971e-010, 9.78221e-010, 9.84471e-010, 9.90721e-010, 9.96971e-010, 1.00322e-009,
+ 1.00947e-009, 1.01572e-009, 1.02197e-009, 1.02822e-009, 1.03447e-009, 1.04072e-009,
+ 1.04697e-009, 1.05322e-009, 1.05947e-009, 1.06572e-009, 1.07197e-009, 1.07822e-009,
+ 1.08447e-009, 1.09072e-009, 1.09697e-009, 1.10322e-009, 1.10947e-009, 1.11572e-009,
+ 1.12197e-009, 1.12822e-009, 1.13447e-009, 1.14072e-009, 1.14697e-009, 1.15322e-009,
+ 1.15947e-009, 1.16572e-009, 1.17197e-009, 1.17822e-009, 1.18447e-009, 1.19072e-009,
+ 1.19697e-009, 1.20322e-009, 1.20947e-009, 1.21572e-009, 1.22197e-009, 1.22822e-009,
+ 1.23447e-009, 1.24072e-009, 1.24697e-009, 1.25322e-009, 1.25947e-009, 1.26572e-009,
+ 1.27197e-009, 1.27822e-009, 1.28447e-009, 1.29072e-009, 1.29697e-009, 1.30322e-009,
+ 1.30947e-009, 1.31572e-009, 1.32197e-009, 1.32822e-009)"
+          kdata_0to1_min="(0, 0.00144844, 0.00161591, 0.00178283, 0.00194921, 0.00211506,
+ 0.0087038, 0.00937234, 0.0100361, 0.0106951, 0.0113493, 0.0221732,
+ 0.0235462, 0.0248913, 0.0262091, 0.027512, 0.0384896, 0.040387,
+ 0.0422566, 0.0440992, 0.0459152, 0.0477052, 0.0909226, 0.0947716,
+ 0.0985008, 0.102115, 0.10562, 0.151672, 0.156561, 0.161263,
+ 0.165788, 0.170143, 0.231451, 0.237879, 0.244041, 0.249991,
+ 0.255738, 0.306646, 0.314487, 0.322133, 0.329544, 0.346723,
+ 0.354268, 0.361647, 0.368849, 0.375871, 0.436727, 0.446473,
+ 0.456075, 0.465528, 0.47489, 0.508024, 0.518296, 0.528421,
+ 0.538431, 0.548284, 0.578952, 0.589365, 0.599555, 0.609511,
+ 0.619187, 0.661993, 0.673295, 0.684356, 0.695153, 0.695174,
+ 0.703634, 0.711667, 0.719248, 0.725866, 0.705895, 0.708557,
+ 0.710598, 0.711564, 0.710588, 0.813801, 0.819259, 0.824199,
+ 0.827163, 0.82912, 0.854347, 0.858385, 0.861996, 0.865003,
+ 0.86646, 0.82184, 0.821897, 0.821674, 0.821592, 0.821429,
+ 0.86842, 0.871631, 0.874676, 0.877554, 0.928498, 0.936229,
+ 0.943903, 0.951517, 0.95907, 0.902802, 0.908617, 0.914903,
+ 0.921194, 0.927466, 0.912617, 0.919099, 0.925592, 0.932094,
+ 0.938605, 0.915914, 0.921739, 0.928803, 0.935927, 0.943095,
+ 0.982139, 0.992066, 1, 1, 0.970056, 0.977633,
+ 0.985279, 0.992996, 1, 0.981505, 0.988024, 0.995008,
+ 1, 1, 0.97652, 0.981778, 0.987072, 0.992403,
+ 0.997772, 0.989569, 0.994141, 0.99874, 1, 1,
+ 0.958503, 0.959695, 0.960888, 0.961952, 0.984313, 0.987439,
+ 0.99058, 0.993734, 0.996902, 0.986424, 0.988754, 0.991091,
+ 0.993435, 0.995786, 0.984205, 0.985709, 0.987216, 0.988726,
+ 0.990238, 0.991754, 0.993272, 0.994792, 0.996316, 0.997843,
+ 0.997771, 0.99948, 1, 1, 0.978729, 0.978557,
+ 0.978385, 0.978213, 0.978042, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 0.984196, 0.983159, 0.982125, 0.981093, 0.980062,
+ 0.991678, 0.991678, 0.991678, 0.991678, 0.991678, 1,
+ 1, 1, 1, 1)"
+          tdata_1to0_min="(1.63161e-011, 2.2246e-011, 2.81759e-011, 3.41058e-011, 4.00356e-011, 4.59655e-011,
+ 5.18954e-011, 5.78253e-011, 6.37551e-011, 6.9685e-011, 7.56149e-011, 8.15448e-011,
+ 8.74746e-011, 9.34045e-011, 9.93344e-011, 1.05264e-010, 1.11194e-010, 1.17124e-010,
+ 1.23054e-010, 1.28984e-010, 1.34914e-010, 1.40843e-010, 1.46773e-010, 1.52703e-010,
+ 1.58633e-010, 1.64563e-010, 1.70493e-010, 1.76423e-010, 1.82353e-010, 1.88282e-010,
+ 1.94212e-010, 2.00142e-010, 2.06072e-010, 2.12002e-010, 2.17932e-010, 2.23862e-010,
+ 2.29792e-010, 2.35721e-010, 2.41651e-010, 2.47581e-010, 2.53511e-010, 2.59441e-010,
+ 2.65371e-010, 2.71301e-010, 2.77231e-010, 2.8316e-010, 2.8909e-010, 2.9502e-010,
+ 3.0095e-010, 3.0688e-010, 3.1281e-010, 3.1874e-010, 3.2467e-010, 3.30599e-010,
+ 3.36529e-010, 3.42459e-010, 3.48389e-010, 3.54319e-010, 3.60249e-010, 3.66179e-010,
+ 3.72109e-010, 3.78038e-010, 3.83968e-010, 3.89898e-010, 3.95828e-010, 4.01758e-010,
+ 4.07688e-010, 4.13618e-010, 4.19548e-010, 4.25477e-010, 4.31407e-010, 4.37337e-010,
+ 4.43267e-010, 4.49197e-010, 4.55127e-010, 4.61057e-010, 4.66987e-010, 4.72916e-010,
+ 4.78846e-010, 4.84776e-010, 4.90706e-010, 4.96636e-010, 5.02566e-010, 5.08496e-010,
+ 5.14426e-010, 5.20355e-010, 5.26285e-010, 5.32215e-010, 5.38145e-010, 5.44075e-010,
+ 5.50005e-010, 5.55935e-010, 5.61865e-010, 5.67794e-010, 5.73724e-010, 5.79654e-010,
+ 5.85584e-010, 5.91514e-010, 5.97444e-010, 6.03374e-010, 6.09304e-010, 6.15233e-010,
+ 6.21163e-010, 6.27093e-010, 6.33023e-010, 6.38953e-010, 6.44883e-010, 6.50813e-010,
+ 6.56743e-010, 6.62672e-010, 6.68602e-010, 6.74532e-010, 6.80462e-010, 6.86392e-010,
+ 6.92322e-010, 6.98252e-010, 7.04182e-010, 7.10111e-010, 7.16041e-010, 7.21971e-010,
+ 7.27901e-010, 7.33831e-010, 7.39761e-010, 7.45691e-010, 7.51621e-010, 7.5755e-010,
+ 7.6348e-010, 7.6941e-010, 7.7534e-010, 7.8127e-010, 7.872e-010, 7.9313e-010,
+ 7.9906e-010, 8.04989e-010, 8.10919e-010, 8.16849e-010, 8.22779e-010, 8.28709e-010,
+ 8.34639e-010, 8.40569e-010, 8.46499e-010, 8.52428e-010, 8.58358e-010, 8.64288e-010,
+ 8.70218e-010, 8.76148e-010, 8.82078e-010, 8.88008e-010, 8.93938e-010, 8.99867e-010,
+ 9.05797e-010, 9.11727e-010, 9.17657e-010, 9.23587e-010, 9.29517e-010, 9.35447e-010,
+ 9.41377e-010, 9.47306e-010, 9.53236e-010, 9.59166e-010, 9.65096e-010, 9.71026e-010,
+ 9.76956e-010, 9.82886e-010, 9.88816e-010, 9.94745e-010, 1.00068e-009, 1.00661e-009,
+ 1.01254e-009, 1.01846e-009, 1.02439e-009, 1.03032e-009, 1.03625e-009, 1.04218e-009,
+ 1.04811e-009, 1.05404e-009, 1.05997e-009, 1.0659e-009, 1.07183e-009, 1.07776e-009,
+ 1.08369e-009, 1.08962e-009, 1.09555e-009, 1.10148e-009, 1.10741e-009, 1.11334e-009,
+ 1.11927e-009, 1.1252e-009, 1.13113e-009, 1.13706e-009, 1.14299e-009, 1.14892e-009,
+ 1.15485e-009, 1.16078e-009, 1.16671e-009, 1.17264e-009, 1.17857e-009, 1.1845e-009,
+ 1.19043e-009, 1.19636e-009, 1.20229e-009, 1.20822e-009)"
+          kdata_1to0_min="(1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 0.944958, 0.941817, 0.939014,
+ 0.936329, 0.933652, 0.928097, 0.926197, 0.924296, 0.922394,
+ 0.920489, 0.918327, 0.916081, 0.742328, 0.734287, 0.726279,
+ 0.718306, 0.710366, 0.5818, 0.572814, 0.563786, 0.554718,
+ 0.545614, 0.432759, 0.422287, 0.411632, 0.400804, 0.390031,
+ 0.357675, 0.345405, 0.33285, 0.319786, 0.306318, 0.299028,
+ 0.281999, 0.263834, 0.245179, 0.224, 0.21373, 0.19043,
+ 0.164822, 0.138767, 0.11283, 0.168453, 0.142421, 0.11653,
+ 0.0898447, 0.064093, 0.12499, 0.101151, 0.0779349, 0.0556811,
+ 0.0329568, 0.116942, 0.0977118, 0.0785584, 0.0587776, 0.0393621,
+ 0.100619, 0.0856291, 0.0698708, 0.0543328, 0.0388455, 0.0738995,
+ 0.0617298, 0.0492707, 0.0366203, 0.0238299, 0.0109021, 0.0561065,
+ 0.0467763, 0.0372812, 0.0274446, 0.0172799, 0.0457196, 0.0381295,
+ 0.0304268, 0.0225745, 0.0145697, 0.0383468, 0.0325389, 0.0266255,
+ 0.0206042, 0.0144643, 0.0365308, 0.0322321, 0.0277894, 0.0232542,
+ 0.0186239, 0.028672, 0.025203, 0.0216809, 0.0181047, 0.0144733,
+ 0.0148853, 0.0116153, 0.00831567, 0.00498609, 0.0016262, 0.0188761,
+ 0.0170186, 0.015139, 0.0132368, 0.0113117, 0.0155086, 0.0140556,
+ 0.0125899, 0.0111111, 0.00961925, 0.0139533, 0.0129102, 0.0118597,
+ 0.0108016, 0.00973602, 0.0114324, 0.0105801, 0.00972376, 0.00886338,
+ 0.00799891, 0.00901914, 0.00830074, 0.00758063, 0.0068588, 0.00613525,
+ 0.00561266, 0.00490209, 0.00419006, 0.00347656, 0.00276158, 0.00173159,
+ 0.000988725, 0.000244458, 0, 0, 0.00391781, 0.00364127,
+ 0.00336415, 0.00308644, 0.00280814, 0.00360153, 0.003408, 0.00321424,
+ 0.00302027, 0.00282607, 0.00282379, 0.00264561, 0.00246717, 0.00228846,
+ 0.00210949, 0.00204093, 0.00187022, 0.00169929, 0.00152814, 0.00135675,
+ 0.00118514, 0.00121595, 0.00106019, 0.000904174, 0.000747895, 0.000591352,
+ 0.00127719, 0.00118284, 0.00108844, 0.000993996, 0.000899505, 0.000727513,
+ 0.000625664, 0.000523821, 0.000421982, 0.000320148, 0.000293503, 0.000198808,
+ 0.000104067, 9.27975e-006, 0, 0.0004531, 0.000407536, 0.000361956,
+ 0.000316359, 0.000270744, 0.000225112, 0)"
+          vdata_min="(-1.8, -1.74, -1.68, -1.62, -1.56, -1.5,
+ -1.44, -1.38, -1.32, -1.26, -1.2, -1.14,
+ -1.08, -1.02, -0.96, -0.9, -0.84, -0.78,
+ -0.72, -0.66, -0.6, -0.54, -0.48, -0.42,
+ -0.36, -0.3, -0.24, -0.18, -0.12, -0.06,
+ 0, 0.06, 0.12, 0.18, 0.24, 0.3,
+ 0.36, 0.42, 0.48, 0.54, 0.6, 0.66,
+ 0.72, 0.78, 0.84, 0.9, 0.96, 1.02,
+ 1.08, 1.14, 1.2, 1.26, 1.32, 1.38,
+ 1.44, 1.5, 1.56, 1.62, 1.68, 1.74,
+ 1.8, 1.86, 1.92, 1.98, 2.04, 2.1,
+ 2.16, 2.22, 2.28, 2.34, 2.4, 2.46,
+ 2.52, 2.58, 2.64, 2.7, 2.76, 2.82,
+ 2.88, 2.94, 3, 3.06, 3.12, 3.18,
+ 3.24, 3.3, 3.36, 3.42, 3.48, 3.54,
+ 3.6)"
+          idata_min="(-2.394, -2.235, -2.075, -1.915, -1.756, -1.596,
+ -1.437, -1.277, -1.118, -0.9586, -0.7993, -0.6403,
+ -0.4841, -0.3375, -0.2096, -0.1333, -0.1135, -0.1032,
+ -0.09427, -0.08574, -0.07761, -0.06996, -0.06286, -0.05631,
+ -0.05017, -0.04422, -0.03837, -0.03258, -0.02687, -0.02127,
+ -0.01578, -0.01053, -0.005574, -0.0009032, 0.003482, 0.007583,
+ 0.0114, 0.01494, 0.0182, 0.02119, 0.0239, 0.02632,
+ 0.02844, 0.03027, 0.03189, 0.03338, 0.03481, 0.0362,
+ 0.03759, 0.03898, 0.04039, 0.04181, 0.04324, 0.0447,
+ 0.04617, 0.04766, 0.04918, 0.05073, 0.0523, 0.0539,
+ 0.05554, 0.05721, 0.05887, 0.06051, 0.06215, 0.06379,
+ 0.06553, 0.06774, 0.07132, 0.07727, 0.08581, 0.09653,
+ 0.109, 0.1233, 0.143, 0.1988, 0.4466, 0.8356,
+ 1.244, 1.664, 2.088, 2.513, 2.938, 3.364,
+ 3.79, 4.216, 4.641, 5.067, 5.493, 5.919,
+ 6.346)"
+          tdata_0to1_max="(7.19709e-011, 7.82209e-011, 8.44709e-011, 9.07209e-011, 9.69709e-011, 1.03221e-010,
+ 1.09471e-010, 1.15721e-010, 1.21971e-010, 1.28221e-010, 1.34471e-010, 1.40721e-010,
+ 1.46971e-010, 1.53221e-010, 1.59471e-010, 1.65721e-010, 1.71971e-010, 1.78221e-010,
+ 1.84471e-010, 1.90721e-010, 1.96971e-010, 2.03221e-010, 2.09471e-010, 2.15721e-010,
+ 2.21971e-010, 2.28221e-010, 2.34471e-010, 2.40721e-010, 2.46971e-010, 2.53221e-010,
+ 2.59471e-010, 2.65721e-010, 2.71971e-010, 2.78221e-010, 2.84471e-010, 2.90721e-010,
+ 2.96971e-010, 3.03221e-010, 3.09471e-010, 3.15721e-010, 3.21971e-010, 3.28221e-010,
+ 3.34471e-010, 3.40721e-010, 3.46971e-010, 3.53221e-010, 3.59471e-010, 3.65721e-010,
+ 3.71971e-010, 3.78221e-010, 3.84471e-010, 3.90721e-010, 3.96971e-010, 4.03221e-010,
+ 4.09471e-010, 4.15721e-010, 4.21971e-010, 4.28221e-010, 4.34471e-010, 4.40721e-010,
+ 4.46971e-010, 4.53221e-010, 4.59471e-010, 4.65721e-010, 4.71971e-010, 4.78221e-010,
+ 4.84471e-010, 4.90721e-010, 4.96971e-010, 5.03221e-010, 5.09471e-010, 5.15721e-010,
+ 5.21971e-010, 5.28221e-010, 5.34471e-010, 5.40721e-010, 5.46971e-010, 5.53221e-010,
+ 5.59471e-010, 5.65721e-010, 5.71971e-010, 5.78221e-010, 5.84471e-010, 5.90721e-010,
+ 5.96971e-010, 6.03221e-010, 6.09471e-010, 6.15721e-010, 6.21971e-010, 6.28221e-010,
+ 6.34471e-010, 6.40721e-010, 6.46971e-010, 6.53221e-010, 6.59471e-010, 6.65721e-010,
+ 6.71971e-010, 6.78221e-010, 6.84471e-010, 6.90721e-010, 6.96971e-010, 7.03221e-010,
+ 7.09471e-010, 7.15721e-010, 7.21971e-010, 7.28221e-010, 7.34471e-010, 7.40721e-010,
+ 7.46971e-010, 7.53221e-010, 7.59471e-010, 7.65721e-010, 7.71971e-010, 7.78221e-010,
+ 7.84471e-010, 7.90721e-010, 7.96971e-010, 8.03221e-010, 8.09471e-010, 8.15721e-010,
+ 8.21971e-010, 8.28221e-010, 8.34471e-010, 8.40721e-010, 8.46971e-010, 8.53221e-010,
+ 8.59471e-010, 8.65721e-010, 8.71971e-010, 8.78221e-010, 8.84471e-010, 8.90721e-010,
+ 8.96971e-010, 9.03221e-010, 9.09471e-010, 9.15721e-010, 9.21971e-010, 9.28221e-010,
+ 9.34471e-010, 9.40721e-010, 9.46971e-010, 9.53221e-010, 9.59471e-010, 9.65721e-010,
+ 9.71971e-010, 9.78221e-010, 9.84471e-010, 9.90721e-010, 9.96971e-010, 1.00322e-009,
+ 1.00947e-009, 1.01572e-009, 1.02197e-009, 1.02822e-009, 1.03447e-009, 1.04072e-009,
+ 1.04697e-009, 1.05322e-009, 1.05947e-009, 1.06572e-009, 1.07197e-009, 1.07822e-009,
+ 1.08447e-009, 1.09072e-009, 1.09697e-009, 1.10322e-009, 1.10947e-009, 1.11572e-009,
+ 1.12197e-009, 1.12822e-009, 1.13447e-009, 1.14072e-009, 1.14697e-009, 1.15322e-009,
+ 1.15947e-009, 1.16572e-009, 1.17197e-009, 1.17822e-009, 1.18447e-009, 1.19072e-009,
+ 1.19697e-009, 1.20322e-009, 1.20947e-009, 1.21572e-009, 1.22197e-009, 1.22822e-009,
+ 1.23447e-009, 1.24072e-009, 1.24697e-009, 1.25322e-009, 1.25947e-009, 1.26572e-009,
+ 1.27197e-009, 1.27822e-009, 1.28447e-009, 1.29072e-009, 1.29697e-009, 1.30322e-009,
+ 1.30947e-009, 1.31572e-009, 1.32197e-009, 1.32822e-009)"
+          kdata_0to1_max="(0, 0.00144844, 0.00161591, 0.00178283, 0.00194921, 0.00211506,
+ 0.0087038, 0.00937234, 0.0100361, 0.0106951, 0.0113493, 0.0221732,
+ 0.0235462, 0.0248913, 0.0262091, 0.027512, 0.0384896, 0.040387,
+ 0.0422566, 0.0440992, 0.0459152, 0.0477052, 0.0909226, 0.0947716,
+ 0.0985008, 0.102115, 0.10562, 0.151672, 0.156561, 0.161263,
+ 0.165788, 0.170143, 0.231451, 0.237879, 0.244041, 0.249991,
+ 0.255738, 0.306646, 0.314487, 0.322133, 0.329544, 0.346723,
+ 0.354268, 0.361647, 0.368849, 0.375871, 0.436727, 0.446473,
+ 0.456075, 0.465528, 0.47489, 0.508024, 0.518296, 0.528421,
+ 0.538431, 0.548284, 0.578952, 0.589365, 0.599555, 0.609511,
+ 0.619187, 0.661993, 0.673295, 0.684356, 0.695153, 0.695174,
+ 0.703634, 0.711667, 0.719248, 0.725866, 0.705895, 0.708557,
+ 0.710598, 0.711564, 0.710588, 0.813801, 0.819259, 0.824199,
+ 0.827163, 0.82912, 0.854347, 0.858385, 0.861996, 0.865003,
+ 0.86646, 0.82184, 0.821897, 0.821674, 0.821592, 0.821429,
+ 0.86842, 0.871631, 0.874676, 0.877554, 0.928498, 0.936229,
+ 0.943903, 0.951517, 0.95907, 0.902802, 0.908617, 0.914903,
+ 0.921194, 0.927466, 0.912617, 0.919099, 0.925592, 0.932094,
+ 0.938605, 0.915914, 0.921739, 0.928803, 0.935927, 0.943095,
+ 0.982139, 0.992066, 1, 1, 0.970056, 0.977633,
+ 0.985279, 0.992996, 1, 0.981505, 0.988024, 0.995008,
+ 1, 1, 0.97652, 0.981778, 0.987072, 0.992403,
+ 0.997772, 0.989569, 0.994141, 0.99874, 1, 1,
+ 0.958503, 0.959695, 0.960888, 0.961952, 0.984313, 0.987439,
+ 0.99058, 0.993734, 0.996902, 0.986424, 0.988754, 0.991091,
+ 0.993435, 0.995786, 0.984205, 0.985709, 0.987216, 0.988726,
+ 0.990238, 0.991754, 0.993272, 0.994792, 0.996316, 0.997843,
+ 0.997771, 0.99948, 1, 1, 0.978729, 0.978557,
+ 0.978385, 0.978213, 0.978042, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 0.984196, 0.983159, 0.982125, 0.981093, 0.980062,
+ 0.991678, 0.991678, 0.991678, 0.991678, 0.991678, 1,
+ 1, 1, 1, 1)"
+          tdata_1to0_max="(1.63161e-011, 2.2246e-011, 2.81759e-011, 3.41058e-011, 4.00356e-011, 4.59655e-011,
+ 5.18954e-011, 5.78253e-011, 6.37551e-011, 6.9685e-011, 7.56149e-011, 8.15448e-011,
+ 8.74746e-011, 9.34045e-011, 9.93344e-011, 1.05264e-010, 1.11194e-010, 1.17124e-010,
+ 1.23054e-010, 1.28984e-010, 1.34914e-010, 1.40843e-010, 1.46773e-010, 1.52703e-010,
+ 1.58633e-010, 1.64563e-010, 1.70493e-010, 1.76423e-010, 1.82353e-010, 1.88282e-010,
+ 1.94212e-010, 2.00142e-010, 2.06072e-010, 2.12002e-010, 2.17932e-010, 2.23862e-010,
+ 2.29792e-010, 2.35721e-010, 2.41651e-010, 2.47581e-010, 2.53511e-010, 2.59441e-010,
+ 2.65371e-010, 2.71301e-010, 2.77231e-010, 2.8316e-010, 2.8909e-010, 2.9502e-010,
+ 3.0095e-010, 3.0688e-010, 3.1281e-010, 3.1874e-010, 3.2467e-010, 3.30599e-010,
+ 3.36529e-010, 3.42459e-010, 3.48389e-010, 3.54319e-010, 3.60249e-010, 3.66179e-010,
+ 3.72109e-010, 3.78038e-010, 3.83968e-010, 3.89898e-010, 3.95828e-010, 4.01758e-010,
+ 4.07688e-010, 4.13618e-010, 4.19548e-010, 4.25477e-010, 4.31407e-010, 4.37337e-010,
+ 4.43267e-010, 4.49197e-010, 4.55127e-010, 4.61057e-010, 4.66987e-010, 4.72916e-010,
+ 4.78846e-010, 4.84776e-010, 4.90706e-010, 4.96636e-010, 5.02566e-010, 5.08496e-010,
+ 5.14426e-010, 5.20355e-010, 5.26285e-010, 5.32215e-010, 5.38145e-010, 5.44075e-010,
+ 5.50005e-010, 5.55935e-010, 5.61865e-010, 5.67794e-010, 5.73724e-010, 5.79654e-010,
+ 5.85584e-010, 5.91514e-010, 5.97444e-010, 6.03374e-010, 6.09304e-010, 6.15233e-010,
+ 6.21163e-010, 6.27093e-010, 6.33023e-010, 6.38953e-010, 6.44883e-010, 6.50813e-010,
+ 6.56743e-010, 6.62672e-010, 6.68602e-010, 6.74532e-010, 6.80462e-010, 6.86392e-010,
+ 6.92322e-010, 6.98252e-010, 7.04182e-010, 7.10111e-010, 7.16041e-010, 7.21971e-010,
+ 7.27901e-010, 7.33831e-010, 7.39761e-010, 7.45691e-010, 7.51621e-010, 7.5755e-010,
+ 7.6348e-010, 7.6941e-010, 7.7534e-010, 7.8127e-010, 7.872e-010, 7.9313e-010,
+ 7.9906e-010, 8.04989e-010, 8.10919e-010, 8.16849e-010, 8.22779e-010, 8.28709e-010,
+ 8.34639e-010, 8.40569e-010, 8.46499e-010, 8.52428e-010, 8.58358e-010, 8.64288e-010,
+ 8.70218e-010, 8.76148e-010, 8.82078e-010, 8.88008e-010, 8.93938e-010, 8.99867e-010,
+ 9.05797e-010, 9.11727e-010, 9.17657e-010, 9.23587e-010, 9.29517e-010, 9.35447e-010,
+ 9.41377e-010, 9.47306e-010, 9.53236e-010, 9.59166e-010, 9.65096e-010, 9.71026e-010,
+ 9.76956e-010, 9.82886e-010, 9.88816e-010, 9.94745e-010, 1.00068e-009, 1.00661e-009,
+ 1.01254e-009, 1.01846e-009, 1.02439e-009, 1.03032e-009, 1.03625e-009, 1.04218e-009,
+ 1.04811e-009, 1.05404e-009, 1.05997e-009, 1.0659e-009, 1.07183e-009, 1.07776e-009,
+ 1.08369e-009, 1.08962e-009, 1.09555e-009, 1.10148e-009, 1.10741e-009, 1.11334e-009,
+ 1.11927e-009, 1.1252e-009, 1.13113e-009, 1.13706e-009, 1.14299e-009, 1.14892e-009,
+ 1.15485e-009, 1.16078e-009, 1.16671e-009, 1.17264e-009, 1.17857e-009, 1.1845e-009,
+ 1.19043e-009, 1.19636e-009, 1.20229e-009, 1.20822e-009)"
+          kdata_1to0_max="(1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 0.944958, 0.941817, 0.939014,
+ 0.936329, 0.933652, 0.928097, 0.926197, 0.924296, 0.922394,
+ 0.920489, 0.918327, 0.916081, 0.742328, 0.734287, 0.726279,
+ 0.718306, 0.710366, 0.5818, 0.572814, 0.563786, 0.554718,
+ 0.545614, 0.432759, 0.422287, 0.411632, 0.400804, 0.390031,
+ 0.357675, 0.345405, 0.33285, 0.319786, 0.306318, 0.299028,
+ 0.281999, 0.263834, 0.245179, 0.224, 0.21373, 0.19043,
+ 0.164822, 0.138767, 0.11283, 0.168453, 0.142421, 0.11653,
+ 0.0898447, 0.064093, 0.12499, 0.101151, 0.0779349, 0.0556811,
+ 0.0329568, 0.116942, 0.0977118, 0.0785584, 0.0587776, 0.0393621,
+ 0.100619, 0.0856291, 0.0698708, 0.0543328, 0.0388455, 0.0738995,
+ 0.0617298, 0.0492707, 0.0366203, 0.0238299, 0.0109021, 0.0561065,
+ 0.0467763, 0.0372812, 0.0274446, 0.0172799, 0.0457196, 0.0381295,
+ 0.0304268, 0.0225745, 0.0145697, 0.0383468, 0.0325389, 0.0266255,
+ 0.0206042, 0.0144643, 0.0365308, 0.0322321, 0.0277894, 0.0232542,
+ 0.0186239, 0.028672, 0.025203, 0.0216809, 0.0181047, 0.0144733,
+ 0.0148853, 0.0116153, 0.00831567, 0.00498609, 0.0016262, 0.0188761,
+ 0.0170186, 0.015139, 0.0132368, 0.0113117, 0.0155086, 0.0140556,
+ 0.0125899, 0.0111111, 0.00961925, 0.0139533, 0.0129102, 0.0118597,
+ 0.0108016, 0.00973602, 0.0114324, 0.0105801, 0.00972376, 0.00886338,
+ 0.00799891, 0.00901914, 0.00830074, 0.00758063, 0.0068588, 0.00613525,
+ 0.00561266, 0.00490209, 0.00419006, 0.00347656, 0.00276158, 0.00173159,
+ 0.000988725, 0.000244458, 0, 0, 0.00391781, 0.00364127,
+ 0.00336415, 0.00308644, 0.00280814, 0.00360153, 0.003408, 0.00321424,
+ 0.00302027, 0.00282607, 0.00282379, 0.00264561, 0.00246717, 0.00228846,
+ 0.00210949, 0.00204093, 0.00187022, 0.00169929, 0.00152814, 0.00135675,
+ 0.00118514, 0.00121595, 0.00106019, 0.000904174, 0.000747895, 0.000591352,
+ 0.00127719, 0.00118284, 0.00108844, 0.000993996, 0.000899505, 0.000727513,
+ 0.000625664, 0.000523821, 0.000421982, 0.000320148, 0.000293503, 0.000198808,
+ 0.000104067, 9.27975e-006, 0, 0.0004531, 0.000407536, 0.000361956,
+ 0.000316359, 0.000270744, 0.000225112, 0)"
+          vdata_max="(-1.8, -1.74, -1.68, -1.62, -1.56, -1.5,
+ -1.44, -1.38, -1.32, -1.26, -1.2, -1.14,
+ -1.08, -1.02, -0.96, -0.9, -0.84, -0.78,
+ -0.72, -0.66, -0.6, -0.54, -0.48, -0.42,
+ -0.36, -0.3, -0.24, -0.18, -0.12, -0.06,
+ 0, 0.06, 0.12, 0.18, 0.24, 0.3,
+ 0.36, 0.42, 0.48, 0.54, 0.6, 0.66,
+ 0.72, 0.78, 0.84, 0.9, 0.96, 1.02,
+ 1.08, 1.14, 1.2, 1.26, 1.32, 1.38,
+ 1.44, 1.5, 1.56, 1.62, 1.68, 1.74,
+ 1.8, 1.86, 1.92, 1.98, 2.04, 2.1,
+ 2.16, 2.22, 2.28, 2.34, 2.4, 2.46,
+ 2.52, 2.58, 2.64, 2.7, 2.76, 2.82,
+ 2.88, 2.94, 3, 3.06, 3.12, 3.18,
+ 3.24, 3.3, 3.36, 3.42, 3.48, 3.54,
+ 3.6)"
+          idata_max="(-2.394, -2.235, -2.075, -1.915, -1.756, -1.596,
+ -1.437, -1.277, -1.118, -0.9586, -0.7993, -0.6403,
+ -0.4841, -0.3375, -0.2096, -0.1333, -0.1135, -0.1032,
+ -0.09427, -0.08574, -0.07761, -0.06996, -0.06286, -0.05631,
+ -0.05017, -0.04422, -0.03837, -0.03258, -0.02687, -0.02127,
+ -0.01578, -0.01053, -0.005574, -0.0009032, 0.003482, 0.007583,
+ 0.0114, 0.01494, 0.0182, 0.02119, 0.0239, 0.02632,
+ 0.02844, 0.03027, 0.03189, 0.03338, 0.03481, 0.0362,
+ 0.03759, 0.03898, 0.04039, 0.04181, 0.04324, 0.0447,
+ 0.04617, 0.04766, 0.04918, 0.05073, 0.0523, 0.0539,
+ 0.05554, 0.05721, 0.05887, 0.06051, 0.06215, 0.06379,
+ 0.06553, 0.06774, 0.07132, 0.07727, 0.08581, 0.09653,
+ 0.109, 0.1233, 0.143, 0.1988, 0.4466, 0.8356,
+ 1.244, 1.664, 2.088, 2.513, 2.938, 3.364,
+ 3.79, 4.216, 4.641, 5.067, 5.493, 5.919,
+ 6.346)"
+ PORT: a_signal
+       a_PuRef
+       d_pullup_control

.model ibis_ktiv(icx_behavioral) MACRO LANG=VHDLAMS LIB=icxbase
.ends MODEL_U6_1

*Define subcircuit for MODEL_U5_1_ip
.subckt MODEL_U5_1_ip a_signal a_control 
VPullUpRef a_PURef 0 1.8
VPullDownRef a_PDRef 0 1e-100


Y_a_control ibis_driver_logic(icx_behavioral)
+ GENERIC: corner="ibis_typ"
+          vmeas_values="( 0.5, 0.5, 0.5 )"
+ PORT: a_control
+       a_gnd
+       d_control

.model ibis_driver_logic(icx_behavioral) MACRO LANG=VHDLAMS LIB=icxbase

X_134 a_signal d_control 0 a_PURef a_PDRef MODEL_U5_1

.ends MODEL_U5_1_ip

*Define subcircuit for MODEL_U5_1
.subckt MODEL_U5_1 a_signal d_control a_gnd a_PURef a_PDRef

C_comp a_signal a_gnd 6e-012

VGCRef a_GCRef 0 0
G_gnd_clamp a_signal a_GCRef table v(a_signal, a_GCRef) = 
+ (-3,0) (1,0) (2,0) 
+ (6,0) 

VPCRef a_PCRef 0 1.8
G_power_clamp a_PCRef a_signal table v(a_PCRef, a_signal) = 
+ (-6,0) (-2,0) (-1,0) 
+ (3,0) 

Y_control ibis_control(icx_behavioral)
+ PORT: d_control
+       d_pullup_control
+       d_pulldown_control

.model ibis_control(icx_behavioral) MACRO LANG=VHDLAMS LIB=icxbase


*IBIS Pulldown tables
Y_PullDown ibis_ktiv(icx_behavioral)
+ GENERIC: corner="ibis_typ"
+          tdata_0to1_typ="(1.63161e-011, 2.2246e-011, 2.81759e-011, 3.41058e-011, 4.00356e-011, 4.59655e-011,
+ 5.18954e-011, 5.78253e-011, 6.37551e-011, 6.9685e-011, 7.56149e-011, 8.15448e-011,
+ 8.74746e-011, 9.34045e-011, 9.93344e-011, 1.05264e-010, 1.11194e-010, 1.17124e-010,
+ 1.23054e-010, 1.28984e-010, 1.34914e-010, 1.40843e-010, 1.46773e-010, 1.52703e-010,
+ 1.58633e-010, 1.64563e-010, 1.70493e-010, 1.76423e-010, 1.82353e-010, 1.88282e-010,
+ 1.94212e-010, 2.00142e-010, 2.06072e-010, 2.12002e-010, 2.17932e-010, 2.23862e-010,
+ 2.29792e-010, 2.35721e-010, 2.41651e-010, 2.47581e-010, 2.53511e-010, 2.59441e-010,
+ 2.65371e-010, 2.71301e-010, 2.77231e-010, 2.8316e-010, 2.8909e-010, 2.9502e-010,
+ 3.0095e-010, 3.0688e-010, 3.1281e-010, 3.1874e-010, 3.2467e-010, 3.30599e-010,
+ 3.36529e-010, 3.42459e-010, 3.48389e-010, 3.54319e-010, 3.60249e-010, 3.66179e-010,
+ 3.72109e-010, 3.78038e-010, 3.83968e-010, 3.89898e-010, 3.95828e-010, 4.01758e-010,
+ 4.07688e-010, 4.13618e-010, 4.19548e-010, 4.25477e-010, 4.31407e-010, 4.37337e-010,
+ 4.43267e-010, 4.49197e-010, 4.55127e-010, 4.61057e-010, 4.66987e-010, 4.72916e-010,
+ 4.78846e-010, 4.84776e-010, 4.90706e-010, 4.96636e-010, 5.02566e-010, 5.08496e-010,
+ 5.14426e-010, 5.20355e-010, 5.26285e-010, 5.32215e-010, 5.38145e-010, 5.44075e-010,
+ 5.50005e-010, 5.55935e-010, 5.61865e-010, 5.67794e-010, 5.73724e-010, 5.79654e-010,
+ 5.85584e-010, 5.91514e-010, 5.97444e-010, 6.03374e-010, 6.09304e-010, 6.15233e-010,
+ 6.21163e-010, 6.27093e-010, 6.33023e-010, 6.38953e-010, 6.44883e-010, 6.50813e-010,
+ 6.56743e-010, 6.62672e-010, 6.68602e-010, 6.74532e-010, 6.80462e-010, 6.86392e-010,
+ 6.92322e-010, 6.98252e-010, 7.04182e-010, 7.10111e-010, 7.16041e-010, 7.21971e-010,
+ 7.27901e-010, 7.33831e-010, 7.39761e-010, 7.45691e-010, 7.51621e-010, 7.5755e-010,
+ 7.6348e-010, 7.6941e-010, 7.7534e-010, 7.8127e-010, 7.872e-010, 7.9313e-010,
+ 7.9906e-010, 8.04989e-010, 8.10919e-010, 8.16849e-010, 8.22779e-010, 8.28709e-010,
+ 8.34639e-010, 8.40569e-010, 8.46499e-010, 8.52428e-010, 8.58358e-010, 8.64288e-010,
+ 8.70218e-010, 8.76148e-010, 8.82078e-010, 8.88008e-010, 8.93938e-010, 8.99867e-010,
+ 9.05797e-010, 9.11727e-010, 9.17657e-010, 9.23587e-010, 9.29517e-010, 9.35447e-010,
+ 9.41377e-010, 9.47306e-010, 9.53236e-010, 9.59166e-010, 9.65096e-010, 9.71026e-010,
+ 9.76956e-010, 9.82886e-010, 9.88816e-010, 9.94745e-010, 1.00068e-009, 1.00661e-009,
+ 1.01254e-009, 1.01846e-009, 1.02439e-009, 1.03032e-009, 1.03625e-009, 1.04218e-009,
+ 1.04811e-009, 1.05404e-009, 1.05997e-009, 1.0659e-009, 1.07183e-009, 1.07776e-009,
+ 1.08369e-009, 1.08962e-009, 1.09555e-009, 1.10148e-009, 1.10741e-009, 1.11334e-009,
+ 1.11927e-009, 1.1252e-009, 1.13113e-009, 1.13706e-009, 1.14299e-009, 1.14892e-009,
+ 1.15485e-009, 1.16078e-009, 1.16671e-009, 1.17264e-009, 1.17857e-009, 1.1845e-009,
+ 1.19043e-009, 1.19636e-009, 1.20229e-009, 1.20822e-009)"
+          kdata_0to1_typ="(0, 0.00693597, 0.00734267, 0.00775038, 0.00815913, 0.00858505,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0.0149774, 0.0168403, 0.0186985, 0.0205519,
+ 0.0224006, 0.0240851, 0.0257124, 0.0534193, 0.0575498, 0.0616171,
+ 0.0656214, 0.069563, 0.102944, 0.109289, 0.1155, 0.121575,
+ 0.127512, 0.185885, 0.194014, 0.201885, 0.209487, 0.216904,
+ 0.262763, 0.270595, 0.278029, 0.284935, 0.291331, 0.389536,
+ 0.397239, 0.403807, 0.409531, 0.41272, 0.458302, 0.460574,
+ 0.460332, 0.45866, 0.456168, 0.521521, 0.519402, 0.516554,
+ 0.512182, 0.507981, 0.562714, 0.560143, 0.557616, 0.556013,
+ 0.55331, 0.659015, 0.662791, 0.666581, 0.669294, 0.672524,
+ 0.716442, 0.724711, 0.731962, 0.740509, 0.749691, 0.739752,
+ 0.749267, 0.759439, 0.770012, 0.780565, 0.791097, 0.79587,
+ 0.809271, 0.822809, 0.836161, 0.849325, 0.834494, 0.847778,
+ 0.862015, 0.876457, 0.891109, 0.864523, 0.877546, 0.890758,
+ 0.904235, 0.918949, 0.917735, 0.932302, 0.946993, 0.961955,
+ 0.977195, 0.924242, 0.935102, 0.946108, 0.957264, 0.968572,
+ 0.909004, 0.915836, 0.922722, 0.929662, 0.936656, 0.952113,
+ 0.960445, 0.968871, 0.977393, 0.986011, 0.960073, 0.966314,
+ 0.972606, 0.97895, 0.985348, 0.970999, 0.976042, 0.98112,
+ 0.986232, 0.991379, 0.972387, 0.975803, 0.979234, 0.98268,
+ 0.986141, 0.967094, 0.968918, 0.970746, 0.972578, 0.974414,
+ 0.973267, 0.97489, 0.976515, 0.978144, 0.979776, 0.98008,
+ 0.981606, 0.983135, 0.984771, 0.986428, 0.984285, 0.985785,
+ 0.987287, 0.988793, 0.990302, 0.982654, 0.983469, 0.984284,
+ 0.9851, 0.985918, 0.989565, 0.990614, 0.991664, 0.992715,
+ 0.993768, 0.993327, 0.994265, 0.995205, 0.996146, 0.997089,
+ 0.998032, 1, 1, 1, 1, 1,
+ 0.99667, 0.997028, 0.997387, 0.997745, 0.998104, 0.993811,
+ 0.993821, 0.99383, 0.99384, 0.993849, 0.998489, 0.998848,
+ 0.999207, 0.999566, 0.999926, 0.998882, 0.999149, 0.999417,
+ 0.999684, 0.999951, 1, 1)"
+          tdata_1to0_typ="(7.19709e-011, 7.82209e-011, 8.44709e-011, 9.07209e-011, 9.69709e-011, 1.03221e-010,
+ 1.09471e-010, 1.15721e-010, 1.21971e-010, 1.28221e-010, 1.34471e-010, 1.40721e-010,
+ 1.46971e-010, 1.53221e-010, 1.59471e-010, 1.65721e-010, 1.71971e-010, 1.78221e-010,
+ 1.84471e-010, 1.90721e-010, 1.96971e-010, 2.03221e-010, 2.09471e-010, 2.15721e-010,
+ 2.21971e-010, 2.28221e-010, 2.34471e-010, 2.40721e-010, 2.46971e-010, 2.53221e-010,
+ 2.59471e-010, 2.65721e-010, 2.71971e-010, 2.78221e-010, 2.84471e-010, 2.90721e-010,
+ 2.96971e-010, 3.03221e-010, 3.09471e-010, 3.15721e-010, 3.21971e-010, 3.28221e-010,
+ 3.34471e-010, 3.40721e-010, 3.46971e-010, 3.53221e-010, 3.59471e-010, 3.65721e-010,
+ 3.71971e-010, 3.78221e-010, 3.84471e-010, 3.90721e-010, 3.96971e-010, 4.03221e-010,
+ 4.09471e-010, 4.15721e-010, 4.21971e-010, 4.28221e-010, 4.34471e-010, 4.40721e-010,
+ 4.46971e-010, 4.53221e-010, 4.59471e-010, 4.65721e-010, 4.71971e-010, 4.78221e-010,
+ 4.84471e-010, 4.90721e-010, 4.96971e-010, 5.03221e-010, 5.09471e-010, 5.15721e-010,
+ 5.21971e-010, 5.28221e-010, 5.34471e-010, 5.40721e-010, 5.46971e-010, 5.53221e-010,
+ 5.59471e-010, 5.65721e-010, 5.71971e-010, 5.78221e-010, 5.84471e-010, 5.90721e-010,
+ 5.96971e-010, 6.03221e-010, 6.09471e-010, 6.15721e-010, 6.21971e-010, 6.28221e-010,
+ 6.34471e-010, 6.40721e-010, 6.46971e-010, 6.53221e-010, 6.59471e-010, 6.65721e-010,
+ 6.71971e-010, 6.78221e-010, 6.84471e-010, 6.90721e-010, 6.96971e-010, 7.03221e-010,
+ 7.09471e-010, 7.15721e-010, 7.21971e-010, 7.28221e-010, 7.34471e-010, 7.40721e-010,
+ 7.46971e-010, 7.53221e-010, 7.59471e-010, 7.65721e-010, 7.71971e-010, 7.78221e-010,
+ 7.84471e-010, 7.90721e-010, 7.96971e-010, 8.03221e-010, 8.09471e-010, 8.15721e-010,
+ 8.21971e-010, 8.28221e-010, 8.34471e-010, 8.40721e-010, 8.46971e-010, 8.53221e-010,
+ 8.59471e-010, 8.65721e-010, 8.71971e-010, 8.78221e-010, 8.84471e-010, 8.90721e-010,
+ 8.96971e-010, 9.03221e-010, 9.09471e-010, 9.15721e-010, 9.21971e-010, 9.28221e-010,
+ 9.34471e-010, 9.40721e-010, 9.46971e-010, 9.53221e-010, 9.59471e-010, 9.65721e-010,
+ 9.71971e-010, 9.78221e-010, 9.84471e-010, 9.90721e-010, 9.96971e-010, 1.00322e-009,
+ 1.00947e-009, 1.01572e-009, 1.02197e-009, 1.02822e-009, 1.03447e-009, 1.04072e-009,
+ 1.04697e-009, 1.05322e-009, 1.05947e-009, 1.06572e-009, 1.07197e-009, 1.07822e-009,
+ 1.08447e-009, 1.09072e-009, 1.09697e-009, 1.10322e-009, 1.10947e-009, 1.11572e-009,
+ 1.12197e-009, 1.12822e-009, 1.13447e-009, 1.14072e-009, 1.14697e-009, 1.15322e-009,
+ 1.15947e-009, 1.16572e-009, 1.17197e-009, 1.17822e-009, 1.18447e-009, 1.19072e-009,
+ 1.19697e-009, 1.20322e-009, 1.20947e-009, 1.21572e-009, 1.22197e-009, 1.22822e-009,
+ 1.23447e-009, 1.24072e-009, 1.24697e-009, 1.25322e-009, 1.25947e-009, 1.26572e-009,
+ 1.27197e-009, 1.27822e-009, 1.28447e-009, 1.29072e-009, 1.29697e-009, 1.30322e-009,
+ 1.30947e-009, 1.31572e-009, 1.32197e-009, 1.32822e-009)"
+          kdata_1to0_typ="(1, 0.969945, 0.967761, 0.965584, 0.963414, 0.961251,
+ 0.922663, 0.917876, 0.913122, 0.908402, 0.903714, 0.851047,
+ 0.843315, 0.835827, 0.828581, 0.821414, 0.777789, 0.768792,
+ 0.759918, 0.751166, 0.742532, 0.734016, 0.55307, 0.537138,
+ 0.52166, 0.506619, 0.491996, 0.366398, 0.350055, 0.334232,
+ 0.318906, 0.304052, 0.267484, 0.253148, 0.23932, 0.225815,
+ 0.212624, 0.239538, 0.228337, 0.217242, 0.206183, 0.204381,
+ 0.194033, 0.183877, 0.173777, 0.163736, 0.198952, 0.190664,
+ 0.182312, 0.1739, 0.165717, 0.170127, 0.16219, 0.154145,
+ 0.146131, 0.138011, 0.141711, 0.13341, 0.124857, 0.116071,
+ 0.107027, 0.153405, 0.145329, 0.136956, 0.128286, 0.11476,
+ 0.103503, 0.0919088, 0.0799865, 0.0670827, 0.0281211, 0.0117597,
+ 0, 0, 0, 0.0834382, 0.0701074, 0.0565091,
+ 0.0408893, 0.0245442, 0.0671925, 0.0543346, 0.0413051, 0.0277456,
+ 0.0127862, 0.00102775, 0, 0, 0, 0,
+ 0.0193647, 0.0104846, 0.00154843, 0, 0.0346995, 0.0293831,
+ 0.0239779, 0.0184849, 0.012905, 0.0133686, 0.00943205, 0.00530731,
+ 0.00108283, 0, 0.00937699, 0.00689617, 0.00437921, 0.00182603,
+ 0, 0.00216168, 0.000431909, 0, 0, 0,
+ 0.0182273, 0.0184874, 0.018742, 0.0189907, 0.0137603, 0.0140486,
+ 0.0143348, 0.014619, 0.0149012, 0.012462, 0.0127637, 0.0131749,
+ 0.0137195, 0.0142671, 0.00858316, 0.00888649, 0.00919061, 0.00949552,
+ 0.00980122, 0.00658873, 0.00668349, 0.00677755, 0.00687091, 0.00696356,
+ 0, 0, 0, 0, 0.0026533, 0.00305218,
+ 0.00345251, 0.00385433, 0.00425764, 0.00128215, 0.00147873, 0.0016757,
+ 0.00187306, 0.00207081, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0.00312929, 0.00354451, 0.00396081, 0.00437819, 0, 0,
+ 0, 0, 0, 0.00283054, 0.00324669, 0.00366393,
+ 0.00408225, 0.00450167, 0.00320158, 0.00351594, 0.00383091, 0.00414651,
+ 0.00446272, 0.00477956, 0.0034087, 0.00361956, 0.0038307, 0.00404212,
+ 0.00425382, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0.00147984,
+ 0.00168904, 0.00189851, 0.00210825, 0)"
+          vdata_typ="(-1.8, -1.74, -1.68, -1.62, -1.56, -1.5,
+ -1.44, -1.38, -1.32, -1.26, -1.2, -1.14,
+ -1.08, -1.02, -0.96, -0.9, -0.84, -0.78,
+ -0.72, -0.66, -0.6, -0.54, -0.48, -0.42,
+ -0.36, -0.3, -0.24, -0.18, -0.12, -0.06,
+ 0, 0.06, 0.12, 0.18, 0.24, 0.3,
+ 0.36, 0.42, 0.48, 0.54, 0.6, 0.66,
+ 0.72, 0.78, 0.84, 0.9, 0.96, 1.02,
+ 1.08, 1.14, 1.2, 1.26, 1.32, 1.38,
+ 1.44, 1.5, 1.56, 1.62, 1.68, 1.74,
+ 1.8, 1.86, 1.92, 1.98, 2.04, 2.1,
+ 2.16, 2.22, 2.28, 2.34, 2.4, 2.46,
+ 2.52, 2.58, 2.64, 2.7, 2.76, 2.82,
+ 2.88, 2.94, 3, 3.06, 3.12, 3.18,
+ 3.24, 3.3, 3.36, 3.42, 3.48, 3.54,
+ 3.6)"
+          idata_typ="(-6.345, -5.918, -5.492, -5.066, -4.64, -4.214,
+ -3.788, -3.363, -2.937, -2.511, -2.086, -1.663,
+ -1.243, -0.8341, -0.4448, -0.196, -0.1389, -0.1177,
+ -0.1018, -0.08764, -0.075, -0.06428, -0.05584, -0.04952,
+ -0.04448, -0.0399, -0.03541, -0.03094, -0.02644, -0.02194,
+ -0.01743, -0.01301, -0.008738, -0.004612, -0.0006315, 0.003204,
+ 0.006895, 0.01044, 0.01383, 0.01707, 0.02014, 0.02303,
+ 0.02573, 0.02821, 0.03045, 0.03244, 0.0342, 0.03576,
+ 0.03718, 0.03853, 0.03986, 0.0412, 0.04257, 0.04398,
+ 0.04543, 0.04695, 0.04854, 0.0502, 0.05195, 0.05377,
+ 0.05569, 0.0577, 0.05975, 0.06183, 0.06393, 0.06606,
+ 0.06826, 0.07067, 0.07359, 0.0773, 0.08184, 0.08709,
+ 0.09294, 0.09942, 0.1074, 0.1257, 0.2032, 0.3338,
+ 0.4821, 0.6392, 0.7982, 0.9575, 1.116, 1.276,
+ 1.435, 1.595, 1.754, 1.914, 2.073, 2.233,
+ 2.392)"
+          tdata_0to1_min="(1.63161e-011, 2.2246e-011, 2.81759e-011, 3.41058e-011, 4.00356e-011, 4.59655e-011,
+ 5.18954e-011, 5.78253e-011, 6.37551e-011, 6.9685e-011, 7.56149e-011, 8.15448e-011,
+ 8.74746e-011, 9.34045e-011, 9.93344e-011, 1.05264e-010, 1.11194e-010, 1.17124e-010,
+ 1.23054e-010, 1.28984e-010, 1.34914e-010, 1.40843e-010, 1.46773e-010, 1.52703e-010,
+ 1.58633e-010, 1.64563e-010, 1.70493e-010, 1.76423e-010, 1.82353e-010, 1.88282e-010,
+ 1.94212e-010, 2.00142e-010, 2.06072e-010, 2.12002e-010, 2.17932e-010, 2.23862e-010,
+ 2.29792e-010, 2.35721e-010, 2.41651e-010, 2.47581e-010, 2.53511e-010, 2.59441e-010,
+ 2.65371e-010, 2.71301e-010, 2.77231e-010, 2.8316e-010, 2.8909e-010, 2.9502e-010,
+ 3.0095e-010, 3.0688e-010, 3.1281e-010, 3.1874e-010, 3.2467e-010, 3.30599e-010,
+ 3.36529e-010, 3.42459e-010, 3.48389e-010, 3.54319e-010, 3.60249e-010, 3.66179e-010,
+ 3.72109e-010, 3.78038e-010, 3.83968e-010, 3.89898e-010, 3.95828e-010, 4.01758e-010,
+ 4.07688e-010, 4.13618e-010, 4.19548e-010, 4.25477e-010, 4.31407e-010, 4.37337e-010,
+ 4.43267e-010, 4.49197e-010, 4.55127e-010, 4.61057e-010, 4.66987e-010, 4.72916e-010,
+ 4.78846e-010, 4.84776e-010, 4.90706e-010, 4.96636e-010, 5.02566e-010, 5.08496e-010,
+ 5.14426e-010, 5.20355e-010, 5.26285e-010, 5.32215e-010, 5.38145e-010, 5.44075e-010,
+ 5.50005e-010, 5.55935e-010, 5.61865e-010, 5.67794e-010, 5.73724e-010, 5.79654e-010,
+ 5.85584e-010, 5.91514e-010, 5.97444e-010, 6.03374e-010, 6.09304e-010, 6.15233e-010,
+ 6.21163e-010, 6.27093e-010, 6.33023e-010, 6.38953e-010, 6.44883e-010, 6.50813e-010,
+ 6.56743e-010, 6.62672e-010, 6.68602e-010, 6.74532e-010, 6.80462e-010, 6.86392e-010,
+ 6.92322e-010, 6.98252e-010, 7.04182e-010, 7.10111e-010, 7.16041e-010, 7.21971e-010,
+ 7.27901e-010, 7.33831e-010, 7.39761e-010, 7.45691e-010, 7.51621e-010, 7.5755e-010,
+ 7.6348e-010, 7.6941e-010, 7.7534e-010, 7.8127e-010, 7.872e-010, 7.9313e-010,
+ 7.9906e-010, 8.04989e-010, 8.10919e-010, 8.16849e-010, 8.22779e-010, 8.28709e-010,
+ 8.34639e-010, 8.40569e-010, 8.46499e-010, 8.52428e-010, 8.58358e-010, 8.64288e-010,
+ 8.70218e-010, 8.76148e-010, 8.82078e-010, 8.88008e-010, 8.93938e-010, 8.99867e-010,
+ 9.05797e-010, 9.11727e-010, 9.17657e-010, 9.23587e-010, 9.29517e-010, 9.35447e-010,
+ 9.41377e-010, 9.47306e-010, 9.53236e-010, 9.59166e-010, 9.65096e-010, 9.71026e-010,
+ 9.76956e-010, 9.82886e-010, 9.88816e-010, 9.94745e-010, 1.00068e-009, 1.00661e-009,
+ 1.01254e-009, 1.01846e-009, 1.02439e-009, 1.03032e-009, 1.03625e-009, 1.04218e-009,
+ 1.04811e-009, 1.05404e-009, 1.05997e-009, 1.0659e-009, 1.07183e-009, 1.07776e-009,
+ 1.08369e-009, 1.08962e-009, 1.09555e-009, 1.10148e-009, 1.10741e-009, 1.11334e-009,
+ 1.11927e-009, 1.1252e-009, 1.13113e-009, 1.13706e-009, 1.14299e-009, 1.14892e-009,
+ 1.15485e-009, 1.16078e-009, 1.16671e-009, 1.17264e-009, 1.17857e-009, 1.1845e-009,
+ 1.19043e-009, 1.19636e-009, 1.20229e-009, 1.20822e-009)"
+          kdata_0to1_min="(0, 0.00693597, 0.00734267, 0.00775038, 0.00815913, 0.00858505,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0.0149774, 0.0168403, 0.0186985, 0.0205519,
+ 0.0224006, 0.0240851, 0.0257124, 0.0534193, 0.0575498, 0.0616171,
+ 0.0656214, 0.069563, 0.102944, 0.109289, 0.1155, 0.121575,
+ 0.127512, 0.185885, 0.194014, 0.201885, 0.209487, 0.216904,
+ 0.262763, 0.270595, 0.278029, 0.284935, 0.291331, 0.389536,
+ 0.397239, 0.403807, 0.409531, 0.41272, 0.458302, 0.460574,
+ 0.460332, 0.45866, 0.456168, 0.521521, 0.519402, 0.516554,
+ 0.512182, 0.507981, 0.562714, 0.560143, 0.557616, 0.556013,
+ 0.55331, 0.659015, 0.662791, 0.666581, 0.669294, 0.672524,
+ 0.716442, 0.724711, 0.731962, 0.740509, 0.749691, 0.739752,
+ 0.749267, 0.759439, 0.770012, 0.780565, 0.791097, 0.79587,
+ 0.809271, 0.822809, 0.836161, 0.849325, 0.834494, 0.847778,
+ 0.862015, 0.876457, 0.891109, 0.864523, 0.877546, 0.890758,
+ 0.904235, 0.918949, 0.917735, 0.932302, 0.946993, 0.961955,
+ 0.977195, 0.924242, 0.935102, 0.946108, 0.957264, 0.968572,
+ 0.909004, 0.915836, 0.922722, 0.929662, 0.936656, 0.952113,
+ 0.960445, 0.968871, 0.977393, 0.986011, 0.960073, 0.966314,
+ 0.972606, 0.97895, 0.985348, 0.970999, 0.976042, 0.98112,
+ 0.986232, 0.991379, 0.972387, 0.975803, 0.979234, 0.98268,
+ 0.986141, 0.967094, 0.968918, 0.970746, 0.972578, 0.974414,
+ 0.973267, 0.97489, 0.976515, 0.978144, 0.979776, 0.98008,
+ 0.981606, 0.983135, 0.984771, 0.986428, 0.984285, 0.985785,
+ 0.987287, 0.988793, 0.990302, 0.982654, 0.983469, 0.984284,
+ 0.9851, 0.985918, 0.989565, 0.990614, 0.991664, 0.992715,
+ 0.993768, 0.993327, 0.994265, 0.995205, 0.996146, 0.997089,
+ 0.998032, 1, 1, 1, 1, 1,
+ 0.99667, 0.997028, 0.997387, 0.997745, 0.998104, 0.993811,
+ 0.993821, 0.99383, 0.99384, 0.993849, 0.998489, 0.998848,
+ 0.999207, 0.999566, 0.999926, 0.998882, 0.999149, 0.999417,
+ 0.999684, 0.999951, 1, 1)"
+          tdata_1to0_min="(7.19709e-011, 7.82209e-011, 8.44709e-011, 9.07209e-011, 9.69709e-011, 1.03221e-010,
+ 1.09471e-010, 1.15721e-010, 1.21971e-010, 1.28221e-010, 1.34471e-010, 1.40721e-010,
+ 1.46971e-010, 1.53221e-010, 1.59471e-010, 1.65721e-010, 1.71971e-010, 1.78221e-010,
+ 1.84471e-010, 1.90721e-010, 1.96971e-010, 2.03221e-010, 2.09471e-010, 2.15721e-010,
+ 2.21971e-010, 2.28221e-010, 2.34471e-010, 2.40721e-010, 2.46971e-010, 2.53221e-010,
+ 2.59471e-010, 2.65721e-010, 2.71971e-010, 2.78221e-010, 2.84471e-010, 2.90721e-010,
+ 2.96971e-010, 3.03221e-010, 3.09471e-010, 3.15721e-010, 3.21971e-010, 3.28221e-010,
+ 3.34471e-010, 3.40721e-010, 3.46971e-010, 3.53221e-010, 3.59471e-010, 3.65721e-010,
+ 3.71971e-010, 3.78221e-010, 3.84471e-010, 3.90721e-010, 3.96971e-010, 4.03221e-010,
+ 4.09471e-010, 4.15721e-010, 4.21971e-010, 4.28221e-010, 4.34471e-010, 4.40721e-010,
+ 4.46971e-010, 4.53221e-010, 4.59471e-010, 4.65721e-010, 4.71971e-010, 4.78221e-010,
+ 4.84471e-010, 4.90721e-010, 4.96971e-010, 5.03221e-010, 5.09471e-010, 5.15721e-010,
+ 5.21971e-010, 5.28221e-010, 5.34471e-010, 5.40721e-010, 5.46971e-010, 5.53221e-010,
+ 5.59471e-010, 5.65721e-010, 5.71971e-010, 5.78221e-010, 5.84471e-010, 5.90721e-010,
+ 5.96971e-010, 6.03221e-010, 6.09471e-010, 6.15721e-010, 6.21971e-010, 6.28221e-010,
+ 6.34471e-010, 6.40721e-010, 6.46971e-010, 6.53221e-010, 6.59471e-010, 6.65721e-010,
+ 6.71971e-010, 6.78221e-010, 6.84471e-010, 6.90721e-010, 6.96971e-010, 7.03221e-010,
+ 7.09471e-010, 7.15721e-010, 7.21971e-010, 7.28221e-010, 7.34471e-010, 7.40721e-010,
+ 7.46971e-010, 7.53221e-010, 7.59471e-010, 7.65721e-010, 7.71971e-010, 7.78221e-010,
+ 7.84471e-010, 7.90721e-010, 7.96971e-010, 8.03221e-010, 8.09471e-010, 8.15721e-010,
+ 8.21971e-010, 8.28221e-010, 8.34471e-010, 8.40721e-010, 8.46971e-010, 8.53221e-010,
+ 8.59471e-010, 8.65721e-010, 8.71971e-010, 8.78221e-010, 8.84471e-010, 8.90721e-010,
+ 8.96971e-010, 9.03221e-010, 9.09471e-010, 9.15721e-010, 9.21971e-010, 9.28221e-010,
+ 9.34471e-010, 9.40721e-010, 9.46971e-010, 9.53221e-010, 9.59471e-010, 9.65721e-010,
+ 9.71971e-010, 9.78221e-010, 9.84471e-010, 9.90721e-010, 9.96971e-010, 1.00322e-009,
+ 1.00947e-009, 1.01572e-009, 1.02197e-009, 1.02822e-009, 1.03447e-009, 1.04072e-009,
+ 1.04697e-009, 1.05322e-009, 1.05947e-009, 1.06572e-009, 1.07197e-009, 1.07822e-009,
+ 1.08447e-009, 1.09072e-009, 1.09697e-009, 1.10322e-009, 1.10947e-009, 1.11572e-009,
+ 1.12197e-009, 1.12822e-009, 1.13447e-009, 1.14072e-009, 1.14697e-009, 1.15322e-009,
+ 1.15947e-009, 1.16572e-009, 1.17197e-009, 1.17822e-009, 1.18447e-009, 1.19072e-009,
+ 1.19697e-009, 1.20322e-009, 1.20947e-009, 1.21572e-009, 1.22197e-009, 1.22822e-009,
+ 1.23447e-009, 1.24072e-009, 1.24697e-009, 1.25322e-009, 1.25947e-009, 1.26572e-009,
+ 1.27197e-009, 1.27822e-009, 1.28447e-009, 1.29072e-009, 1.29697e-009, 1.30322e-009,
+ 1.30947e-009, 1.31572e-009, 1.32197e-009, 1.32822e-009)"
+          kdata_1to0_min="(1, 0.969945, 0.967761, 0.965584, 0.963414, 0.961251,
+ 0.922663, 0.917876, 0.913122, 0.908402, 0.903714, 0.851047,
+ 0.843315, 0.835827, 0.828581, 0.821414, 0.777789, 0.768792,
+ 0.759918, 0.751166, 0.742532, 0.734016, 0.55307, 0.537138,
+ 0.52166, 0.506619, 0.491996, 0.366398, 0.350055, 0.334232,
+ 0.318906, 0.304052, 0.267484, 0.253148, 0.23932, 0.225815,
+ 0.212624, 0.239538, 0.228337, 0.217242, 0.206183, 0.204381,
+ 0.194033, 0.183877, 0.173777, 0.163736, 0.198952, 0.190664,
+ 0.182312, 0.1739, 0.165717, 0.170127, 0.16219, 0.154145,
+ 0.146131, 0.138011, 0.141711, 0.13341, 0.124857, 0.116071,
+ 0.107027, 0.153405, 0.145329, 0.136956, 0.128286, 0.11476,
+ 0.103503, 0.0919088, 0.0799865, 0.0670827, 0.0281211, 0.0117597,
+ 0, 0, 0, 0.0834382, 0.0701074, 0.0565091,
+ 0.0408893, 0.0245442, 0.0671925, 0.0543346, 0.0413051, 0.0277456,
+ 0.0127862, 0.00102775, 0, 0, 0, 0,
+ 0.0193647, 0.0104846, 0.00154843, 0, 0.0346995, 0.0293831,
+ 0.0239779, 0.0184849, 0.012905, 0.0133686, 0.00943205, 0.00530731,
+ 0.00108283, 0, 0.00937699, 0.00689617, 0.00437921, 0.00182603,
+ 0, 0.00216168, 0.000431909, 0, 0, 0,
+ 0.0182273, 0.0184874, 0.018742, 0.0189907, 0.0137603, 0.0140486,
+ 0.0143348, 0.014619, 0.0149012, 0.012462, 0.0127637, 0.0131749,
+ 0.0137195, 0.0142671, 0.00858316, 0.00888649, 0.00919061, 0.00949552,
+ 0.00980122, 0.00658873, 0.00668349, 0.00677755, 0.00687091, 0.00696356,
+ 0, 0, 0, 0, 0.0026533, 0.00305218,
+ 0.00345251, 0.00385433, 0.00425764, 0.00128215, 0.00147873, 0.0016757,
+ 0.00187306, 0.00207081, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0.00312929, 0.00354451, 0.00396081, 0.00437819, 0, 0,
+ 0, 0, 0, 0.00283054, 0.00324669, 0.00366393,
+ 0.00408225, 0.00450167, 0.00320158, 0.00351594, 0.00383091, 0.00414651,
+ 0.00446272, 0.00477956, 0.0034087, 0.00361956, 0.0038307, 0.00404212,
+ 0.00425382, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0.00147984,
+ 0.00168904, 0.00189851, 0.00210825, 0)"
+          vdata_min="(-1.8, -1.74, -1.68, -1.62, -1.56, -1.5,
+ -1.44, -1.38, -1.32, -1.26, -1.2, -1.14,
+ -1.08, -1.02, -0.96, -0.9, -0.84, -0.78,
+ -0.72, -0.66, -0.6, -0.54, -0.48, -0.42,
+ -0.36, -0.3, -0.24, -0.18, -0.12, -0.06,
+ 0, 0.06, 0.12, 0.18, 0.24, 0.3,
+ 0.36, 0.42, 0.48, 0.54, 0.6, 0.66,
+ 0.72, 0.78, 0.84, 0.9, 0.96, 1.02,
+ 1.08, 1.14, 1.2, 1.26, 1.32, 1.38,
+ 1.44, 1.5, 1.56, 1.62, 1.68, 1.74,
+ 1.8, 1.86, 1.92, 1.98, 2.04, 2.1,
+ 2.16, 2.22, 2.28, 2.34, 2.4, 2.46,
+ 2.52, 2.58, 2.64, 2.7, 2.76, 2.82,
+ 2.88, 2.94, 3, 3.06, 3.12, 3.18,
+ 3.24, 3.3, 3.36, 3.42, 3.48, 3.54,
+ 3.6)"
+          idata_min="(-6.345, -5.918, -5.492, -5.066, -4.64, -4.214,
+ -3.788, -3.363, -2.937, -2.511, -2.086, -1.663,
+ -1.243, -0.8341, -0.4448, -0.196, -0.1389, -0.1177,
+ -0.1018, -0.08764, -0.075, -0.06428, -0.05584, -0.04952,
+ -0.04448, -0.0399, -0.03541, -0.03094, -0.02644, -0.02194,
+ -0.01743, -0.01301, -0.008738, -0.004612, -0.0006315, 0.003204,
+ 0.006895, 0.01044, 0.01383, 0.01707, 0.02014, 0.02303,
+ 0.02573, 0.02821, 0.03045, 0.03244, 0.0342, 0.03576,
+ 0.03718, 0.03853, 0.03986, 0.0412, 0.04257, 0.04398,
+ 0.04543, 0.04695, 0.04854, 0.0502, 0.05195, 0.05377,
+ 0.05569, 0.0577, 0.05975, 0.06183, 0.06393, 0.06606,
+ 0.06826, 0.07067, 0.07359, 0.0773, 0.08184, 0.08709,
+ 0.09294, 0.09942, 0.1074, 0.1257, 0.2032, 0.3338,
+ 0.4821, 0.6392, 0.7982, 0.9575, 1.116, 1.276,
+ 1.435, 1.595, 1.754, 1.914, 2.073, 2.233,
+ 2.392)"
+          tdata_0to1_max="(1.63161e-011, 2.2246e-011, 2.81759e-011, 3.41058e-011, 4.00356e-011, 4.59655e-011,
+ 5.18954e-011, 5.78253e-011, 6.37551e-011, 6.9685e-011, 7.56149e-011, 8.15448e-011,
+ 8.74746e-011, 9.34045e-011, 9.93344e-011, 1.05264e-010, 1.11194e-010, 1.17124e-010,
+ 1.23054e-010, 1.28984e-010, 1.34914e-010, 1.40843e-010, 1.46773e-010, 1.52703e-010,
+ 1.58633e-010, 1.64563e-010, 1.70493e-010, 1.76423e-010, 1.82353e-010, 1.88282e-010,
+ 1.94212e-010, 2.00142e-010, 2.06072e-010, 2.12002e-010, 2.17932e-010, 2.23862e-010,
+ 2.29792e-010, 2.35721e-010, 2.41651e-010, 2.47581e-010, 2.53511e-010, 2.59441e-010,
+ 2.65371e-010, 2.71301e-010, 2.77231e-010, 2.8316e-010, 2.8909e-010, 2.9502e-010,
+ 3.0095e-010, 3.0688e-010, 3.1281e-010, 3.1874e-010, 3.2467e-010, 3.30599e-010,
+ 3.36529e-010, 3.42459e-010, 3.48389e-010, 3.54319e-010, 3.60249e-010, 3.66179e-010,
+ 3.72109e-010, 3.78038e-010, 3.83968e-010, 3.89898e-010, 3.95828e-010, 4.01758e-010,
+ 4.07688e-010, 4.13618e-010, 4.19548e-010, 4.25477e-010, 4.31407e-010, 4.37337e-010,
+ 4.43267e-010, 4.49197e-010, 4.55127e-010, 4.61057e-010, 4.66987e-010, 4.72916e-010,
+ 4.78846e-010, 4.84776e-010, 4.90706e-010, 4.96636e-010, 5.02566e-010, 5.08496e-010,
+ 5.14426e-010, 5.20355e-010, 5.26285e-010, 5.32215e-010, 5.38145e-010, 5.44075e-010,
+ 5.50005e-010, 5.55935e-010, 5.61865e-010, 5.67794e-010, 5.73724e-010, 5.79654e-010,
+ 5.85584e-010, 5.91514e-010, 5.97444e-010, 6.03374e-010, 6.09304e-010, 6.15233e-010,
+ 6.21163e-010, 6.27093e-010, 6.33023e-010, 6.38953e-010, 6.44883e-010, 6.50813e-010,
+ 6.56743e-010, 6.62672e-010, 6.68602e-010, 6.74532e-010, 6.80462e-010, 6.86392e-010,
+ 6.92322e-010, 6.98252e-010, 7.04182e-010, 7.10111e-010, 7.16041e-010, 7.21971e-010,
+ 7.27901e-010, 7.33831e-010, 7.39761e-010, 7.45691e-010, 7.51621e-010, 7.5755e-010,
+ 7.6348e-010, 7.6941e-010, 7.7534e-010, 7.8127e-010, 7.872e-010, 7.9313e-010,
+ 7.9906e-010, 8.04989e-010, 8.10919e-010, 8.16849e-010, 8.22779e-010, 8.28709e-010,
+ 8.34639e-010, 8.40569e-010, 8.46499e-010, 8.52428e-010, 8.58358e-010, 8.64288e-010,
+ 8.70218e-010, 8.76148e-010, 8.82078e-010, 8.88008e-010, 8.93938e-010, 8.99867e-010,
+ 9.05797e-010, 9.11727e-010, 9.17657e-010, 9.23587e-010, 9.29517e-010, 9.35447e-010,
+ 9.41377e-010, 9.47306e-010, 9.53236e-010, 9.59166e-010, 9.65096e-010, 9.71026e-010,
+ 9.76956e-010, 9.82886e-010, 9.88816e-010, 9.94745e-010, 1.00068e-009, 1.00661e-009,
+ 1.01254e-009, 1.01846e-009, 1.02439e-009, 1.03032e-009, 1.03625e-009, 1.04218e-009,
+ 1.04811e-009, 1.05404e-009, 1.05997e-009, 1.0659e-009, 1.07183e-009, 1.07776e-009,
+ 1.08369e-009, 1.08962e-009, 1.09555e-009, 1.10148e-009, 1.10741e-009, 1.11334e-009,
+ 1.11927e-009, 1.1252e-009, 1.13113e-009, 1.13706e-009, 1.14299e-009, 1.14892e-009,
+ 1.15485e-009, 1.16078e-009, 1.16671e-009, 1.17264e-009, 1.17857e-009, 1.1845e-009,
+ 1.19043e-009, 1.19636e-009, 1.20229e-009, 1.20822e-009)"
+          kdata_0to1_max="(0, 0.00693597, 0.00734267, 0.00775038, 0.00815913, 0.00858505,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0.0149774, 0.0168403, 0.0186985, 0.0205519,
+ 0.0224006, 0.0240851, 0.0257124, 0.0534193, 0.0575498, 0.0616171,
+ 0.0656214, 0.069563, 0.102944, 0.109289, 0.1155, 0.121575,
+ 0.127512, 0.185885, 0.194014, 0.201885, 0.209487, 0.216904,
+ 0.262763, 0.270595, 0.278029, 0.284935, 0.291331, 0.389536,
+ 0.397239, 0.403807, 0.409531, 0.41272, 0.458302, 0.460574,
+ 0.460332, 0.45866, 0.456168, 0.521521, 0.519402, 0.516554,
+ 0.512182, 0.507981, 0.562714, 0.560143, 0.557616, 0.556013,
+ 0.55331, 0.659015, 0.662791, 0.666581, 0.669294, 0.672524,
+ 0.716442, 0.724711, 0.731962, 0.740509, 0.749691, 0.739752,
+ 0.749267, 0.759439, 0.770012, 0.780565, 0.791097, 0.79587,
+ 0.809271, 0.822809, 0.836161, 0.849325, 0.834494, 0.847778,
+ 0.862015, 0.876457, 0.891109, 0.864523, 0.877546, 0.890758,
+ 0.904235, 0.918949, 0.917735, 0.932302, 0.946993, 0.961955,
+ 0.977195, 0.924242, 0.935102, 0.946108, 0.957264, 0.968572,
+ 0.909004, 0.915836, 0.922722, 0.929662, 0.936656, 0.952113,
+ 0.960445, 0.968871, 0.977393, 0.986011, 0.960073, 0.966314,
+ 0.972606, 0.97895, 0.985348, 0.970999, 0.976042, 0.98112,
+ 0.986232, 0.991379, 0.972387, 0.975803, 0.979234, 0.98268,
+ 0.986141, 0.967094, 0.968918, 0.970746, 0.972578, 0.974414,
+ 0.973267, 0.97489, 0.976515, 0.978144, 0.979776, 0.98008,
+ 0.981606, 0.983135, 0.984771, 0.986428, 0.984285, 0.985785,
+ 0.987287, 0.988793, 0.990302, 0.982654, 0.983469, 0.984284,
+ 0.9851, 0.985918, 0.989565, 0.990614, 0.991664, 0.992715,
+ 0.993768, 0.993327, 0.994265, 0.995205, 0.996146, 0.997089,
+ 0.998032, 1, 1, 1, 1, 1,
+ 0.99667, 0.997028, 0.997387, 0.997745, 0.998104, 0.993811,
+ 0.993821, 0.99383, 0.99384, 0.993849, 0.998489, 0.998848,
+ 0.999207, 0.999566, 0.999926, 0.998882, 0.999149, 0.999417,
+ 0.999684, 0.999951, 1, 1)"
+          tdata_1to0_max="(7.19709e-011, 7.82209e-011, 8.44709e-011, 9.07209e-011, 9.69709e-011, 1.03221e-010,
+ 1.09471e-010, 1.15721e-010, 1.21971e-010, 1.28221e-010, 1.34471e-010, 1.40721e-010,
+ 1.46971e-010, 1.53221e-010, 1.59471e-010, 1.65721e-010, 1.71971e-010, 1.78221e-010,
+ 1.84471e-010, 1.90721e-010, 1.96971e-010, 2.03221e-010, 2.09471e-010, 2.15721e-010,
+ 2.21971e-010, 2.28221e-010, 2.34471e-010, 2.40721e-010, 2.46971e-010, 2.53221e-010,
+ 2.59471e-010, 2.65721e-010, 2.71971e-010, 2.78221e-010, 2.84471e-010, 2.90721e-010,
+ 2.96971e-010, 3.03221e-010, 3.09471e-010, 3.15721e-010, 3.21971e-010, 3.28221e-010,
+ 3.34471e-010, 3.40721e-010, 3.46971e-010, 3.53221e-010, 3.59471e-010, 3.65721e-010,
+ 3.71971e-010, 3.78221e-010, 3.84471e-010, 3.90721e-010, 3.96971e-010, 4.03221e-010,
+ 4.09471e-010, 4.15721e-010, 4.21971e-010, 4.28221e-010, 4.34471e-010, 4.40721e-010,
+ 4.46971e-010, 4.53221e-010, 4.59471e-010, 4.65721e-010, 4.71971e-010, 4.78221e-010,
+ 4.84471e-010, 4.90721e-010, 4.96971e-010, 5.03221e-010, 5.09471e-010, 5.15721e-010,
+ 5.21971e-010, 5.28221e-010, 5.34471e-010, 5.40721e-010, 5.46971e-010, 5.53221e-010,
+ 5.59471e-010, 5.65721e-010, 5.71971e-010, 5.78221e-010, 5.84471e-010, 5.90721e-010,
+ 5.96971e-010, 6.03221e-010, 6.09471e-010, 6.15721e-010, 6.21971e-010, 6.28221e-010,
+ 6.34471e-010, 6.40721e-010, 6.46971e-010, 6.53221e-010, 6.59471e-010, 6.65721e-010,
+ 6.71971e-010, 6.78221e-010, 6.84471e-010, 6.90721e-010, 6.96971e-010, 7.03221e-010,
+ 7.09471e-010, 7.15721e-010, 7.21971e-010, 7.28221e-010, 7.34471e-010, 7.40721e-010,
+ 7.46971e-010, 7.53221e-010, 7.59471e-010, 7.65721e-010, 7.71971e-010, 7.78221e-010,
+ 7.84471e-010, 7.90721e-010, 7.96971e-010, 8.03221e-010, 8.09471e-010, 8.15721e-010,
+ 8.21971e-010, 8.28221e-010, 8.34471e-010, 8.40721e-010, 8.46971e-010, 8.53221e-010,
+ 8.59471e-010, 8.65721e-010, 8.71971e-010, 8.78221e-010, 8.84471e-010, 8.90721e-010,
+ 8.96971e-010, 9.03221e-010, 9.09471e-010, 9.15721e-010, 9.21971e-010, 9.28221e-010,
+ 9.34471e-010, 9.40721e-010, 9.46971e-010, 9.53221e-010, 9.59471e-010, 9.65721e-010,
+ 9.71971e-010, 9.78221e-010, 9.84471e-010, 9.90721e-010, 9.96971e-010, 1.00322e-009,
+ 1.00947e-009, 1.01572e-009, 1.02197e-009, 1.02822e-009, 1.03447e-009, 1.04072e-009,
+ 1.04697e-009, 1.05322e-009, 1.05947e-009, 1.06572e-009, 1.07197e-009, 1.07822e-009,
+ 1.08447e-009, 1.09072e-009, 1.09697e-009, 1.10322e-009, 1.10947e-009, 1.11572e-009,
+ 1.12197e-009, 1.12822e-009, 1.13447e-009, 1.14072e-009, 1.14697e-009, 1.15322e-009,
+ 1.15947e-009, 1.16572e-009, 1.17197e-009, 1.17822e-009, 1.18447e-009, 1.19072e-009,
+ 1.19697e-009, 1.20322e-009, 1.20947e-009, 1.21572e-009, 1.22197e-009, 1.22822e-009,
+ 1.23447e-009, 1.24072e-009, 1.24697e-009, 1.25322e-009, 1.25947e-009, 1.26572e-009,
+ 1.27197e-009, 1.27822e-009, 1.28447e-009, 1.29072e-009, 1.29697e-009, 1.30322e-009,
+ 1.30947e-009, 1.31572e-009, 1.32197e-009, 1.32822e-009)"
+          kdata_1to0_max="(1, 0.969945, 0.967761, 0.965584, 0.963414, 0.961251,
+ 0.922663, 0.917876, 0.913122, 0.908402, 0.903714, 0.851047,
+ 0.843315, 0.835827, 0.828581, 0.821414, 0.777789, 0.768792,
+ 0.759918, 0.751166, 0.742532, 0.734016, 0.55307, 0.537138,
+ 0.52166, 0.506619, 0.491996, 0.366398, 0.350055, 0.334232,
+ 0.318906, 0.304052, 0.267484, 0.253148, 0.23932, 0.225815,
+ 0.212624, 0.239538, 0.228337, 0.217242, 0.206183, 0.204381,
+ 0.194033, 0.183877, 0.173777, 0.163736, 0.198952, 0.190664,
+ 0.182312, 0.1739, 0.165717, 0.170127, 0.16219, 0.154145,
+ 0.146131, 0.138011, 0.141711, 0.13341, 0.124857, 0.116071,
+ 0.107027, 0.153405, 0.145329, 0.136956, 0.128286, 0.11476,
+ 0.103503, 0.0919088, 0.0799865, 0.0670827, 0.0281211, 0.0117597,
+ 0, 0, 0, 0.0834382, 0.0701074, 0.0565091,
+ 0.0408893, 0.0245442, 0.0671925, 0.0543346, 0.0413051, 0.0277456,
+ 0.0127862, 0.00102775, 0, 0, 0, 0,
+ 0.0193647, 0.0104846, 0.00154843, 0, 0.0346995, 0.0293831,
+ 0.0239779, 0.0184849, 0.012905, 0.0133686, 0.00943205, 0.00530731,
+ 0.00108283, 0, 0.00937699, 0.00689617, 0.00437921, 0.00182603,
+ 0, 0.00216168, 0.000431909, 0, 0, 0,
+ 0.0182273, 0.0184874, 0.018742, 0.0189907, 0.0137603, 0.0140486,
+ 0.0143348, 0.014619, 0.0149012, 0.012462, 0.0127637, 0.0131749,
+ 0.0137195, 0.0142671, 0.00858316, 0.00888649, 0.00919061, 0.00949552,
+ 0.00980122, 0.00658873, 0.00668349, 0.00677755, 0.00687091, 0.00696356,
+ 0, 0, 0, 0, 0.0026533, 0.00305218,
+ 0.00345251, 0.00385433, 0.00425764, 0.00128215, 0.00147873, 0.0016757,
+ 0.00187306, 0.00207081, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0.00312929, 0.00354451, 0.00396081, 0.00437819, 0, 0,
+ 0, 0, 0, 0.00283054, 0.00324669, 0.00366393,
+ 0.00408225, 0.00450167, 0.00320158, 0.00351594, 0.00383091, 0.00414651,
+ 0.00446272, 0.00477956, 0.0034087, 0.00361956, 0.0038307, 0.00404212,
+ 0.00425382, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0.00147984,
+ 0.00168904, 0.00189851, 0.00210825, 0)"
+          vdata_max="(-1.8, -1.74, -1.68, -1.62, -1.56, -1.5,
+ -1.44, -1.38, -1.32, -1.26, -1.2, -1.14,
+ -1.08, -1.02, -0.96, -0.9, -0.84, -0.78,
+ -0.72, -0.66, -0.6, -0.54, -0.48, -0.42,
+ -0.36, -0.3, -0.24, -0.18, -0.12, -0.06,
+ 0, 0.06, 0.12, 0.18, 0.24, 0.3,
+ 0.36, 0.42, 0.48, 0.54, 0.6, 0.66,
+ 0.72, 0.78, 0.84, 0.9, 0.96, 1.02,
+ 1.08, 1.14, 1.2, 1.26, 1.32, 1.38,
+ 1.44, 1.5, 1.56, 1.62, 1.68, 1.74,
+ 1.8, 1.86, 1.92, 1.98, 2.04, 2.1,
+ 2.16, 2.22, 2.28, 2.34, 2.4, 2.46,
+ 2.52, 2.58, 2.64, 2.7, 2.76, 2.82,
+ 2.88, 2.94, 3, 3.06, 3.12, 3.18,
+ 3.24, 3.3, 3.36, 3.42, 3.48, 3.54,
+ 3.6)"
+          idata_max="(-6.345, -5.918, -5.492, -5.066, -4.64, -4.214,
+ -3.788, -3.363, -2.937, -2.511, -2.086, -1.663,
+ -1.243, -0.8341, -0.4448, -0.196, -0.1389, -0.1177,
+ -0.1018, -0.08764, -0.075, -0.06428, -0.05584, -0.04952,
+ -0.04448, -0.0399, -0.03541, -0.03094, -0.02644, -0.02194,
+ -0.01743, -0.01301, -0.008738, -0.004612, -0.0006315, 0.003204,
+ 0.006895, 0.01044, 0.01383, 0.01707, 0.02014, 0.02303,
+ 0.02573, 0.02821, 0.03045, 0.03244, 0.0342, 0.03576,
+ 0.03718, 0.03853, 0.03986, 0.0412, 0.04257, 0.04398,
+ 0.04543, 0.04695, 0.04854, 0.0502, 0.05195, 0.05377,
+ 0.05569, 0.0577, 0.05975, 0.06183, 0.06393, 0.06606,
+ 0.06826, 0.07067, 0.07359, 0.0773, 0.08184, 0.08709,
+ 0.09294, 0.09942, 0.1074, 0.1257, 0.2032, 0.3338,
+ 0.4821, 0.6392, 0.7982, 0.9575, 1.116, 1.276,
+ 1.435, 1.595, 1.754, 1.914, 2.073, 2.233,
+ 2.392)"
+ PORT: a_PdRef
+       a_signal
+       d_pulldown_control


*IBIS Pullup tables
Y_PullUp ibis_ktiv(icx_behavioral)
+ GENERIC: corner="ibis_typ"
+          tdata_0to1_typ="(7.19709e-011, 7.82209e-011, 8.44709e-011, 9.07209e-011, 9.69709e-011, 1.03221e-010,
+ 1.09471e-010, 1.15721e-010, 1.21971e-010, 1.28221e-010, 1.34471e-010, 1.40721e-010,
+ 1.46971e-010, 1.53221e-010, 1.59471e-010, 1.65721e-010, 1.71971e-010, 1.78221e-010,
+ 1.84471e-010, 1.90721e-010, 1.96971e-010, 2.03221e-010, 2.09471e-010, 2.15721e-010,
+ 2.21971e-010, 2.28221e-010, 2.34471e-010, 2.40721e-010, 2.46971e-010, 2.53221e-010,
+ 2.59471e-010, 2.65721e-010, 2.71971e-010, 2.78221e-010, 2.84471e-010, 2.90721e-010,
+ 2.96971e-010, 3.03221e-010, 3.09471e-010, 3.15721e-010, 3.21971e-010, 3.28221e-010,
+ 3.34471e-010, 3.40721e-010, 3.46971e-010, 3.53221e-010, 3.59471e-010, 3.65721e-010,
+ 3.71971e-010, 3.78221e-010, 3.84471e-010, 3.90721e-010, 3.96971e-010, 4.03221e-010,
+ 4.09471e-010, 4.15721e-010, 4.21971e-010, 4.28221e-010, 4.34471e-010, 4.40721e-010,
+ 4.46971e-010, 4.53221e-010, 4.59471e-010, 4.65721e-010, 4.71971e-010, 4.78221e-010,
+ 4.84471e-010, 4.90721e-010, 4.96971e-010, 5.03221e-010, 5.09471e-010, 5.15721e-010,
+ 5.21971e-010, 5.28221e-010, 5.34471e-010, 5.40721e-010, 5.46971e-010, 5.53221e-010,
+ 5.59471e-010, 5.65721e-010, 5.71971e-010, 5.78221e-010, 5.84471e-010, 5.90721e-010,
+ 5.96971e-010, 6.03221e-010, 6.09471e-010, 6.15721e-010, 6.21971e-010, 6.28221e-010,
+ 6.34471e-010, 6.40721e-010, 6.46971e-010, 6.53221e-010, 6.59471e-010, 6.65721e-010,
+ 6.71971e-010, 6.78221e-010, 6.84471e-010, 6.90721e-010, 6.96971e-010, 7.03221e-010,
+ 7.09471e-010, 7.15721e-010, 7.21971e-010, 7.28221e-010, 7.34471e-010, 7.40721e-010,
+ 7.46971e-010, 7.53221e-010, 7.59471e-010, 7.65721e-010, 7.71971e-010, 7.78221e-010,
+ 7.84471e-010, 7.90721e-010, 7.96971e-010, 8.03221e-010, 8.09471e-010, 8.15721e-010,
+ 8.21971e-010, 8.28221e-010, 8.34471e-010, 8.40721e-010, 8.46971e-010, 8.53221e-010,
+ 8.59471e-010, 8.65721e-010, 8.71971e-010, 8.78221e-010, 8.84471e-010, 8.90721e-010,
+ 8.96971e-010, 9.03221e-010, 9.09471e-010, 9.15721e-010, 9.21971e-010, 9.28221e-010,
+ 9.34471e-010, 9.40721e-010, 9.46971e-010, 9.53221e-010, 9.59471e-010, 9.65721e-010,
+ 9.71971e-010, 9.78221e-010, 9.84471e-010, 9.90721e-010, 9.96971e-010, 1.00322e-009,
+ 1.00947e-009, 1.01572e-009, 1.02197e-009, 1.02822e-009, 1.03447e-009, 1.04072e-009,
+ 1.04697e-009, 1.05322e-009, 1.05947e-009, 1.06572e-009, 1.07197e-009, 1.07822e-009,
+ 1.08447e-009, 1.09072e-009, 1.09697e-009, 1.10322e-009, 1.10947e-009, 1.11572e-009,
+ 1.12197e-009, 1.12822e-009, 1.13447e-009, 1.14072e-009, 1.14697e-009, 1.15322e-009,
+ 1.15947e-009, 1.16572e-009, 1.17197e-009, 1.17822e-009, 1.18447e-009, 1.19072e-009,
+ 1.19697e-009, 1.20322e-009, 1.20947e-009, 1.21572e-009, 1.22197e-009, 1.22822e-009,
+ 1.23447e-009, 1.24072e-009, 1.24697e-009, 1.25322e-009, 1.25947e-009, 1.26572e-009,
+ 1.27197e-009, 1.27822e-009, 1.28447e-009, 1.29072e-009, 1.29697e-009, 1.30322e-009,
+ 1.30947e-009, 1.31572e-009, 1.32197e-009, 1.32822e-009)"
+          kdata_0to1_typ="(0, 0.00144844, 0.00161591, 0.00178283, 0.00194921, 0.00211506,
+ 0.0087038, 0.00937234, 0.0100361, 0.0106951, 0.0113493, 0.0221732,
+ 0.0235462, 0.0248913, 0.0262091, 0.027512, 0.0384896, 0.040387,
+ 0.0422566, 0.0440992, 0.0459152, 0.0477052, 0.0909226, 0.0947716,
+ 0.0985008, 0.102115, 0.10562, 0.151672, 0.156561, 0.161263,
+ 0.165788, 0.170143, 0.231451, 0.237879, 0.244041, 0.249991,
+ 0.255738, 0.306646, 0.314487, 0.322133, 0.329544, 0.346723,
+ 0.354268, 0.361647, 0.368849, 0.375871, 0.436727, 0.446473,
+ 0.456075, 0.465528, 0.47489, 0.508024, 0.518296, 0.528421,
+ 0.538431, 0.548284, 0.578952, 0.589365, 0.599555, 0.609511,
+ 0.619187, 0.661993, 0.673295, 0.684356, 0.695153, 0.695174,
+ 0.703634, 0.711667, 0.719248, 0.725866, 0.705895, 0.708557,
+ 0.710598, 0.711564, 0.710588, 0.813801, 0.819259, 0.824199,
+ 0.827163, 0.82912, 0.854347, 0.858385, 0.861996, 0.865003,
+ 0.86646, 0.82184, 0.821897, 0.821674, 0.821592, 0.821429,
+ 0.86842, 0.871631, 0.874676, 0.877554, 0.928498, 0.936229,
+ 0.943903, 0.951517, 0.95907, 0.902802, 0.908617, 0.914903,
+ 0.921194, 0.927466, 0.912617, 0.919099, 0.925592, 0.932094,
+ 0.938605, 0.915914, 0.921739, 0.928803, 0.935927, 0.943095,
+ 0.982139, 0.992066, 1, 1, 0.970056, 0.977633,
+ 0.985279, 0.992996, 1, 0.981505, 0.988024, 0.995008,
+ 1, 1, 0.97652, 0.981778, 0.987072, 0.992403,
+ 0.997772, 0.989569, 0.994141, 0.99874, 1, 1,
+ 0.958503, 0.959695, 0.960888, 0.961952, 0.984313, 0.987439,
+ 0.99058, 0.993734, 0.996902, 0.986424, 0.988754, 0.991091,
+ 0.993435, 0.995786, 0.984205, 0.985709, 0.987216, 0.988726,
+ 0.990238, 0.991754, 0.993272, 0.994792, 0.996316, 0.997843,
+ 0.997771, 0.99948, 1, 1, 0.978729, 0.978557,
+ 0.978385, 0.978213, 0.978042, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 0.984196, 0.983159, 0.982125, 0.981093, 0.980062,
+ 0.991678, 0.991678, 0.991678, 0.991678, 0.991678, 1,
+ 1, 1, 1, 1)"
+          tdata_1to0_typ="(1.63161e-011, 2.2246e-011, 2.81759e-011, 3.41058e-011, 4.00356e-011, 4.59655e-011,
+ 5.18954e-011, 5.78253e-011, 6.37551e-011, 6.9685e-011, 7.56149e-011, 8.15448e-011,
+ 8.74746e-011, 9.34045e-011, 9.93344e-011, 1.05264e-010, 1.11194e-010, 1.17124e-010,
+ 1.23054e-010, 1.28984e-010, 1.34914e-010, 1.40843e-010, 1.46773e-010, 1.52703e-010,
+ 1.58633e-010, 1.64563e-010, 1.70493e-010, 1.76423e-010, 1.82353e-010, 1.88282e-010,
+ 1.94212e-010, 2.00142e-010, 2.06072e-010, 2.12002e-010, 2.17932e-010, 2.23862e-010,
+ 2.29792e-010, 2.35721e-010, 2.41651e-010, 2.47581e-010, 2.53511e-010, 2.59441e-010,
+ 2.65371e-010, 2.71301e-010, 2.77231e-010, 2.8316e-010, 2.8909e-010, 2.9502e-010,
+ 3.0095e-010, 3.0688e-010, 3.1281e-010, 3.1874e-010, 3.2467e-010, 3.30599e-010,
+ 3.36529e-010, 3.42459e-010, 3.48389e-010, 3.54319e-010, 3.60249e-010, 3.66179e-010,
+ 3.72109e-010, 3.78038e-010, 3.83968e-010, 3.89898e-010, 3.95828e-010, 4.01758e-010,
+ 4.07688e-010, 4.13618e-010, 4.19548e-010, 4.25477e-010, 4.31407e-010, 4.37337e-010,
+ 4.43267e-010, 4.49197e-010, 4.55127e-010, 4.61057e-010, 4.66987e-010, 4.72916e-010,
+ 4.78846e-010, 4.84776e-010, 4.90706e-010, 4.96636e-010, 5.02566e-010, 5.08496e-010,
+ 5.14426e-010, 5.20355e-010, 5.26285e-010, 5.32215e-010, 5.38145e-010, 5.44075e-010,
+ 5.50005e-010, 5.55935e-010, 5.61865e-010, 5.67794e-010, 5.73724e-010, 5.79654e-010,
+ 5.85584e-010, 5.91514e-010, 5.97444e-010, 6.03374e-010, 6.09304e-010, 6.15233e-010,
+ 6.21163e-010, 6.27093e-010, 6.33023e-010, 6.38953e-010, 6.44883e-010, 6.50813e-010,
+ 6.56743e-010, 6.62672e-010, 6.68602e-010, 6.74532e-010, 6.80462e-010, 6.86392e-010,
+ 6.92322e-010, 6.98252e-010, 7.04182e-010, 7.10111e-010, 7.16041e-010, 7.21971e-010,
+ 7.27901e-010, 7.33831e-010, 7.39761e-010, 7.45691e-010, 7.51621e-010, 7.5755e-010,
+ 7.6348e-010, 7.6941e-010, 7.7534e-010, 7.8127e-010, 7.872e-010, 7.9313e-010,
+ 7.9906e-010, 8.04989e-010, 8.10919e-010, 8.16849e-010, 8.22779e-010, 8.28709e-010,
+ 8.34639e-010, 8.40569e-010, 8.46499e-010, 8.52428e-010, 8.58358e-010, 8.64288e-010,
+ 8.70218e-010, 8.76148e-010, 8.82078e-010, 8.88008e-010, 8.93938e-010, 8.99867e-010,
+ 9.05797e-010, 9.11727e-010, 9.17657e-010, 9.23587e-010, 9.29517e-010, 9.35447e-010,
+ 9.41377e-010, 9.47306e-010, 9.53236e-010, 9.59166e-010, 9.65096e-010, 9.71026e-010,
+ 9.76956e-010, 9.82886e-010, 9.88816e-010, 9.94745e-010, 1.00068e-009, 1.00661e-009,
+ 1.01254e-009, 1.01846e-009, 1.02439e-009, 1.03032e-009, 1.03625e-009, 1.04218e-009,
+ 1.04811e-009, 1.05404e-009, 1.05997e-009, 1.0659e-009, 1.07183e-009, 1.07776e-009,
+ 1.08369e-009, 1.08962e-009, 1.09555e-009, 1.10148e-009, 1.10741e-009, 1.11334e-009,
+ 1.11927e-009, 1.1252e-009, 1.13113e-009, 1.13706e-009, 1.14299e-009, 1.14892e-009,
+ 1.15485e-009, 1.16078e-009, 1.16671e-009, 1.17264e-009, 1.17857e-009, 1.1845e-009,
+ 1.19043e-009, 1.19636e-009, 1.20229e-009, 1.20822e-009)"
+          kdata_1to0_typ="(1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 0.944958, 0.941817, 0.939014,
+ 0.936329, 0.933652, 0.928097, 0.926197, 0.924296, 0.922394,
+ 0.920489, 0.918327, 0.916081, 0.742328, 0.734287, 0.726279,
+ 0.718306, 0.710366, 0.5818, 0.572814, 0.563786, 0.554718,
+ 0.545614, 0.432759, 0.422287, 0.411632, 0.400804, 0.390031,
+ 0.357675, 0.345405, 0.33285, 0.319786, 0.306318, 0.299028,
+ 0.281999, 0.263834, 0.245179, 0.224, 0.21373, 0.19043,
+ 0.164822, 0.138767, 0.11283, 0.168453, 0.142421, 0.11653,
+ 0.0898447, 0.064093, 0.12499, 0.101151, 0.0779349, 0.0556811,
+ 0.0329568, 0.116942, 0.0977118, 0.0785584, 0.0587776, 0.0393621,
+ 0.100619, 0.0856291, 0.0698708, 0.0543328, 0.0388455, 0.0738995,
+ 0.0617298, 0.0492707, 0.0366203, 0.0238299, 0.0109021, 0.0561065,
+ 0.0467763, 0.0372812, 0.0274446, 0.0172799, 0.0457196, 0.0381295,
+ 0.0304268, 0.0225745, 0.0145697, 0.0383468, 0.0325389, 0.0266255,
+ 0.0206042, 0.0144643, 0.0365308, 0.0322321, 0.0277894, 0.0232542,
+ 0.0186239, 0.028672, 0.025203, 0.0216809, 0.0181047, 0.0144733,
+ 0.0148853, 0.0116153, 0.00831567, 0.00498609, 0.0016262, 0.0188761,
+ 0.0170186, 0.015139, 0.0132368, 0.0113117, 0.0155086, 0.0140556,
+ 0.0125899, 0.0111111, 0.00961925, 0.0139533, 0.0129102, 0.0118597,
+ 0.0108016, 0.00973602, 0.0114324, 0.0105801, 0.00972376, 0.00886338,
+ 0.00799891, 0.00901914, 0.00830074, 0.00758063, 0.0068588, 0.00613525,
+ 0.00561266, 0.00490209, 0.00419006, 0.00347656, 0.00276158, 0.00173159,
+ 0.000988725, 0.000244458, 0, 0, 0.00391781, 0.00364127,
+ 0.00336415, 0.00308644, 0.00280814, 0.00360153, 0.003408, 0.00321424,
+ 0.00302027, 0.00282607, 0.00282379, 0.00264561, 0.00246717, 0.00228846,
+ 0.00210949, 0.00204093, 0.00187022, 0.00169929, 0.00152814, 0.00135675,
+ 0.00118514, 0.00121595, 0.00106019, 0.000904174, 0.000747895, 0.000591352,
+ 0.00127719, 0.00118284, 0.00108844, 0.000993996, 0.000899505, 0.000727513,
+ 0.000625664, 0.000523821, 0.000421982, 0.000320148, 0.000293503, 0.000198808,
+ 0.000104067, 9.27975e-006, 0, 0.0004531, 0.000407536, 0.000361956,
+ 0.000316359, 0.000270744, 0.000225112, 0)"
+          vdata_typ="(-1.8, -1.74, -1.68, -1.62, -1.56, -1.5,
+ -1.44, -1.38, -1.32, -1.26, -1.2, -1.14,
+ -1.08, -1.02, -0.96, -0.9, -0.84, -0.78,
+ -0.72, -0.66, -0.6, -0.54, -0.48, -0.42,
+ -0.36, -0.3, -0.24, -0.18, -0.12, -0.06,
+ 0, 0.06, 0.12, 0.18, 0.24, 0.3,
+ 0.36, 0.42, 0.48, 0.54, 0.6, 0.66,
+ 0.72, 0.78, 0.84, 0.9, 0.96, 1.02,
+ 1.08, 1.14, 1.2, 1.26, 1.32, 1.38,
+ 1.44, 1.5, 1.56, 1.62, 1.68, 1.74,
+ 1.8, 1.86, 1.92, 1.98, 2.04, 2.1,
+ 2.16, 2.22, 2.28, 2.34, 2.4, 2.46,
+ 2.52, 2.58, 2.64, 2.7, 2.76, 2.82,
+ 2.88, 2.94, 3, 3.06, 3.12, 3.18,
+ 3.24, 3.3, 3.36, 3.42, 3.48, 3.54,
+ 3.6)"
+          idata_typ="(-2.394, -2.235, -2.075, -1.915, -1.756, -1.596,
+ -1.437, -1.277, -1.118, -0.9586, -0.7993, -0.6403,
+ -0.4841, -0.3375, -0.2096, -0.1333, -0.1135, -0.1032,
+ -0.09427, -0.08574, -0.07761, -0.06996, -0.06286, -0.05631,
+ -0.05017, -0.04422, -0.03837, -0.03258, -0.02687, -0.02127,
+ -0.01578, -0.01053, -0.005574, -0.0009032, 0.003482, 0.007583,
+ 0.0114, 0.01494, 0.0182, 0.02119, 0.0239, 0.02632,
+ 0.02844, 0.03027, 0.03189, 0.03338, 0.03481, 0.0362,
+ 0.03759, 0.03898, 0.04039, 0.04181, 0.04324, 0.0447,
+ 0.04617, 0.04766, 0.04918, 0.05073, 0.0523, 0.0539,
+ 0.05554, 0.05721, 0.05887, 0.06051, 0.06215, 0.06379,
+ 0.06553, 0.06774, 0.07132, 0.07727, 0.08581, 0.09653,
+ 0.109, 0.1233, 0.143, 0.1988, 0.4466, 0.8356,
+ 1.244, 1.664, 2.088, 2.513, 2.938, 3.364,
+ 3.79, 4.216, 4.641, 5.067, 5.493, 5.919,
+ 6.346)"
+          tdata_0to1_min="(7.19709e-011, 7.82209e-011, 8.44709e-011, 9.07209e-011, 9.69709e-011, 1.03221e-010,
+ 1.09471e-010, 1.15721e-010, 1.21971e-010, 1.28221e-010, 1.34471e-010, 1.40721e-010,
+ 1.46971e-010, 1.53221e-010, 1.59471e-010, 1.65721e-010, 1.71971e-010, 1.78221e-010,
+ 1.84471e-010, 1.90721e-010, 1.96971e-010, 2.03221e-010, 2.09471e-010, 2.15721e-010,
+ 2.21971e-010, 2.28221e-010, 2.34471e-010, 2.40721e-010, 2.46971e-010, 2.53221e-010,
+ 2.59471e-010, 2.65721e-010, 2.71971e-010, 2.78221e-010, 2.84471e-010, 2.90721e-010,
+ 2.96971e-010, 3.03221e-010, 3.09471e-010, 3.15721e-010, 3.21971e-010, 3.28221e-010,
+ 3.34471e-010, 3.40721e-010, 3.46971e-010, 3.53221e-010, 3.59471e-010, 3.65721e-010,
+ 3.71971e-010, 3.78221e-010, 3.84471e-010, 3.90721e-010, 3.96971e-010, 4.03221e-010,
+ 4.09471e-010, 4.15721e-010, 4.21971e-010, 4.28221e-010, 4.34471e-010, 4.40721e-010,
+ 4.46971e-010, 4.53221e-010, 4.59471e-010, 4.65721e-010, 4.71971e-010, 4.78221e-010,
+ 4.84471e-010, 4.90721e-010, 4.96971e-010, 5.03221e-010, 5.09471e-010, 5.15721e-010,
+ 5.21971e-010, 5.28221e-010, 5.34471e-010, 5.40721e-010, 5.46971e-010, 5.53221e-010,
+ 5.59471e-010, 5.65721e-010, 5.71971e-010, 5.78221e-010, 5.84471e-010, 5.90721e-010,
+ 5.96971e-010, 6.03221e-010, 6.09471e-010, 6.15721e-010, 6.21971e-010, 6.28221e-010,
+ 6.34471e-010, 6.40721e-010, 6.46971e-010, 6.53221e-010, 6.59471e-010, 6.65721e-010,
+ 6.71971e-010, 6.78221e-010, 6.84471e-010, 6.90721e-010, 6.96971e-010, 7.03221e-010,
+ 7.09471e-010, 7.15721e-010, 7.21971e-010, 7.28221e-010, 7.34471e-010, 7.40721e-010,
+ 7.46971e-010, 7.53221e-010, 7.59471e-010, 7.65721e-010, 7.71971e-010, 7.78221e-010,
+ 7.84471e-010, 7.90721e-010, 7.96971e-010, 8.03221e-010, 8.09471e-010, 8.15721e-010,
+ 8.21971e-010, 8.28221e-010, 8.34471e-010, 8.40721e-010, 8.46971e-010, 8.53221e-010,
+ 8.59471e-010, 8.65721e-010, 8.71971e-010, 8.78221e-010, 8.84471e-010, 8.90721e-010,
+ 8.96971e-010, 9.03221e-010, 9.09471e-010, 9.15721e-010, 9.21971e-010, 9.28221e-010,
+ 9.34471e-010, 9.40721e-010, 9.46971e-010, 9.53221e-010, 9.59471e-010, 9.65721e-010,
+ 9.71971e-010, 9.78221e-010, 9.84471e-010, 9.90721e-010, 9.96971e-010, 1.00322e-009,
+ 1.00947e-009, 1.01572e-009, 1.02197e-009, 1.02822e-009, 1.03447e-009, 1.04072e-009,
+ 1.04697e-009, 1.05322e-009, 1.05947e-009, 1.06572e-009, 1.07197e-009, 1.07822e-009,
+ 1.08447e-009, 1.09072e-009, 1.09697e-009, 1.10322e-009, 1.10947e-009, 1.11572e-009,
+ 1.12197e-009, 1.12822e-009, 1.13447e-009, 1.14072e-009, 1.14697e-009, 1.15322e-009,
+ 1.15947e-009, 1.16572e-009, 1.17197e-009, 1.17822e-009, 1.18447e-009, 1.19072e-009,
+ 1.19697e-009, 1.20322e-009, 1.20947e-009, 1.21572e-009, 1.22197e-009, 1.22822e-009,
+ 1.23447e-009, 1.24072e-009, 1.24697e-009, 1.25322e-009, 1.25947e-009, 1.26572e-009,
+ 1.27197e-009, 1.27822e-009, 1.28447e-009, 1.29072e-009, 1.29697e-009, 1.30322e-009,
+ 1.30947e-009, 1.31572e-009, 1.32197e-009, 1.32822e-009)"
+          kdata_0to1_min="(0, 0.00144844, 0.00161591, 0.00178283, 0.00194921, 0.00211506,
+ 0.0087038, 0.00937234, 0.0100361, 0.0106951, 0.0113493, 0.0221732,
+ 0.0235462, 0.0248913, 0.0262091, 0.027512, 0.0384896, 0.040387,
+ 0.0422566, 0.0440992, 0.0459152, 0.0477052, 0.0909226, 0.0947716,
+ 0.0985008, 0.102115, 0.10562, 0.151672, 0.156561, 0.161263,
+ 0.165788, 0.170143, 0.231451, 0.237879, 0.244041, 0.249991,
+ 0.255738, 0.306646, 0.314487, 0.322133, 0.329544, 0.346723,
+ 0.354268, 0.361647, 0.368849, 0.375871, 0.436727, 0.446473,
+ 0.456075, 0.465528, 0.47489, 0.508024, 0.518296, 0.528421,
+ 0.538431, 0.548284, 0.578952, 0.589365, 0.599555, 0.609511,
+ 0.619187, 0.661993, 0.673295, 0.684356, 0.695153, 0.695174,
+ 0.703634, 0.711667, 0.719248, 0.725866, 0.705895, 0.708557,
+ 0.710598, 0.711564, 0.710588, 0.813801, 0.819259, 0.824199,
+ 0.827163, 0.82912, 0.854347, 0.858385, 0.861996, 0.865003,
+ 0.86646, 0.82184, 0.821897, 0.821674, 0.821592, 0.821429,
+ 0.86842, 0.871631, 0.874676, 0.877554, 0.928498, 0.936229,
+ 0.943903, 0.951517, 0.95907, 0.902802, 0.908617, 0.914903,
+ 0.921194, 0.927466, 0.912617, 0.919099, 0.925592, 0.932094,
+ 0.938605, 0.915914, 0.921739, 0.928803, 0.935927, 0.943095,
+ 0.982139, 0.992066, 1, 1, 0.970056, 0.977633,
+ 0.985279, 0.992996, 1, 0.981505, 0.988024, 0.995008,
+ 1, 1, 0.97652, 0.981778, 0.987072, 0.992403,
+ 0.997772, 0.989569, 0.994141, 0.99874, 1, 1,
+ 0.958503, 0.959695, 0.960888, 0.961952, 0.984313, 0.987439,
+ 0.99058, 0.993734, 0.996902, 0.986424, 0.988754, 0.991091,
+ 0.993435, 0.995786, 0.984205, 0.985709, 0.987216, 0.988726,
+ 0.990238, 0.991754, 0.993272, 0.994792, 0.996316, 0.997843,
+ 0.997771, 0.99948, 1, 1, 0.978729, 0.978557,
+ 0.978385, 0.978213, 0.978042, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 0.984196, 0.983159, 0.982125, 0.981093, 0.980062,
+ 0.991678, 0.991678, 0.991678, 0.991678, 0.991678, 1,
+ 1, 1, 1, 1)"
+          tdata_1to0_min="(1.63161e-011, 2.2246e-011, 2.81759e-011, 3.41058e-011, 4.00356e-011, 4.59655e-011,
+ 5.18954e-011, 5.78253e-011, 6.37551e-011, 6.9685e-011, 7.56149e-011, 8.15448e-011,
+ 8.74746e-011, 9.34045e-011, 9.93344e-011, 1.05264e-010, 1.11194e-010, 1.17124e-010,
+ 1.23054e-010, 1.28984e-010, 1.34914e-010, 1.40843e-010, 1.46773e-010, 1.52703e-010,
+ 1.58633e-010, 1.64563e-010, 1.70493e-010, 1.76423e-010, 1.82353e-010, 1.88282e-010,
+ 1.94212e-010, 2.00142e-010, 2.06072e-010, 2.12002e-010, 2.17932e-010, 2.23862e-010,
+ 2.29792e-010, 2.35721e-010, 2.41651e-010, 2.47581e-010, 2.53511e-010, 2.59441e-010,
+ 2.65371e-010, 2.71301e-010, 2.77231e-010, 2.8316e-010, 2.8909e-010, 2.9502e-010,
+ 3.0095e-010, 3.0688e-010, 3.1281e-010, 3.1874e-010, 3.2467e-010, 3.30599e-010,
+ 3.36529e-010, 3.42459e-010, 3.48389e-010, 3.54319e-010, 3.60249e-010, 3.66179e-010,
+ 3.72109e-010, 3.78038e-010, 3.83968e-010, 3.89898e-010, 3.95828e-010, 4.01758e-010,
+ 4.07688e-010, 4.13618e-010, 4.19548e-010, 4.25477e-010, 4.31407e-010, 4.37337e-010,
+ 4.43267e-010, 4.49197e-010, 4.55127e-010, 4.61057e-010, 4.66987e-010, 4.72916e-010,
+ 4.78846e-010, 4.84776e-010, 4.90706e-010, 4.96636e-010, 5.02566e-010, 5.08496e-010,
+ 5.14426e-010, 5.20355e-010, 5.26285e-010, 5.32215e-010, 5.38145e-010, 5.44075e-010,
+ 5.50005e-010, 5.55935e-010, 5.61865e-010, 5.67794e-010, 5.73724e-010, 5.79654e-010,
+ 5.85584e-010, 5.91514e-010, 5.97444e-010, 6.03374e-010, 6.09304e-010, 6.15233e-010,
+ 6.21163e-010, 6.27093e-010, 6.33023e-010, 6.38953e-010, 6.44883e-010, 6.50813e-010,
+ 6.56743e-010, 6.62672e-010, 6.68602e-010, 6.74532e-010, 6.80462e-010, 6.86392e-010,
+ 6.92322e-010, 6.98252e-010, 7.04182e-010, 7.10111e-010, 7.16041e-010, 7.21971e-010,
+ 7.27901e-010, 7.33831e-010, 7.39761e-010, 7.45691e-010, 7.51621e-010, 7.5755e-010,
+ 7.6348e-010, 7.6941e-010, 7.7534e-010, 7.8127e-010, 7.872e-010, 7.9313e-010,
+ 7.9906e-010, 8.04989e-010, 8.10919e-010, 8.16849e-010, 8.22779e-010, 8.28709e-010,
+ 8.34639e-010, 8.40569e-010, 8.46499e-010, 8.52428e-010, 8.58358e-010, 8.64288e-010,
+ 8.70218e-010, 8.76148e-010, 8.82078e-010, 8.88008e-010, 8.93938e-010, 8.99867e-010,
+ 9.05797e-010, 9.11727e-010, 9.17657e-010, 9.23587e-010, 9.29517e-010, 9.35447e-010,
+ 9.41377e-010, 9.47306e-010, 9.53236e-010, 9.59166e-010, 9.65096e-010, 9.71026e-010,
+ 9.76956e-010, 9.82886e-010, 9.88816e-010, 9.94745e-010, 1.00068e-009, 1.00661e-009,
+ 1.01254e-009, 1.01846e-009, 1.02439e-009, 1.03032e-009, 1.03625e-009, 1.04218e-009,
+ 1.04811e-009, 1.05404e-009, 1.05997e-009, 1.0659e-009, 1.07183e-009, 1.07776e-009,
+ 1.08369e-009, 1.08962e-009, 1.09555e-009, 1.10148e-009, 1.10741e-009, 1.11334e-009,
+ 1.11927e-009, 1.1252e-009, 1.13113e-009, 1.13706e-009, 1.14299e-009, 1.14892e-009,
+ 1.15485e-009, 1.16078e-009, 1.16671e-009, 1.17264e-009, 1.17857e-009, 1.1845e-009,
+ 1.19043e-009, 1.19636e-009, 1.20229e-009, 1.20822e-009)"
+          kdata_1to0_min="(1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 0.944958, 0.941817, 0.939014,
+ 0.936329, 0.933652, 0.928097, 0.926197, 0.924296, 0.922394,
+ 0.920489, 0.918327, 0.916081, 0.742328, 0.734287, 0.726279,
+ 0.718306, 0.710366, 0.5818, 0.572814, 0.563786, 0.554718,
+ 0.545614, 0.432759, 0.422287, 0.411632, 0.400804, 0.390031,
+ 0.357675, 0.345405, 0.33285, 0.319786, 0.306318, 0.299028,
+ 0.281999, 0.263834, 0.245179, 0.224, 0.21373, 0.19043,
+ 0.164822, 0.138767, 0.11283, 0.168453, 0.142421, 0.11653,
+ 0.0898447, 0.064093, 0.12499, 0.101151, 0.0779349, 0.0556811,
+ 0.0329568, 0.116942, 0.0977118, 0.0785584, 0.0587776, 0.0393621,
+ 0.100619, 0.0856291, 0.0698708, 0.0543328, 0.0388455, 0.0738995,
+ 0.0617298, 0.0492707, 0.0366203, 0.0238299, 0.0109021, 0.0561065,
+ 0.0467763, 0.0372812, 0.0274446, 0.0172799, 0.0457196, 0.0381295,
+ 0.0304268, 0.0225745, 0.0145697, 0.0383468, 0.0325389, 0.0266255,
+ 0.0206042, 0.0144643, 0.0365308, 0.0322321, 0.0277894, 0.0232542,
+ 0.0186239, 0.028672, 0.025203, 0.0216809, 0.0181047, 0.0144733,
+ 0.0148853, 0.0116153, 0.00831567, 0.00498609, 0.0016262, 0.0188761,
+ 0.0170186, 0.015139, 0.0132368, 0.0113117, 0.0155086, 0.0140556,
+ 0.0125899, 0.0111111, 0.00961925, 0.0139533, 0.0129102, 0.0118597,
+ 0.0108016, 0.00973602, 0.0114324, 0.0105801, 0.00972376, 0.00886338,
+ 0.00799891, 0.00901914, 0.00830074, 0.00758063, 0.0068588, 0.00613525,
+ 0.00561266, 0.00490209, 0.00419006, 0.00347656, 0.00276158, 0.00173159,
+ 0.000988725, 0.000244458, 0, 0, 0.00391781, 0.00364127,
+ 0.00336415, 0.00308644, 0.00280814, 0.00360153, 0.003408, 0.00321424,
+ 0.00302027, 0.00282607, 0.00282379, 0.00264561, 0.00246717, 0.00228846,
+ 0.00210949, 0.00204093, 0.00187022, 0.00169929, 0.00152814, 0.00135675,
+ 0.00118514, 0.00121595, 0.00106019, 0.000904174, 0.000747895, 0.000591352,
+ 0.00127719, 0.00118284, 0.00108844, 0.000993996, 0.000899505, 0.000727513,
+ 0.000625664, 0.000523821, 0.000421982, 0.000320148, 0.000293503, 0.000198808,
+ 0.000104067, 9.27975e-006, 0, 0.0004531, 0.000407536, 0.000361956,
+ 0.000316359, 0.000270744, 0.000225112, 0)"
+          vdata_min="(-1.8, -1.74, -1.68, -1.62, -1.56, -1.5,
+ -1.44, -1.38, -1.32, -1.26, -1.2, -1.14,
+ -1.08, -1.02, -0.96, -0.9, -0.84, -0.78,
+ -0.72, -0.66, -0.6, -0.54, -0.48, -0.42,
+ -0.36, -0.3, -0.24, -0.18, -0.12, -0.06,
+ 0, 0.06, 0.12, 0.18, 0.24, 0.3,
+ 0.36, 0.42, 0.48, 0.54, 0.6, 0.66,
+ 0.72, 0.78, 0.84, 0.9, 0.96, 1.02,
+ 1.08, 1.14, 1.2, 1.26, 1.32, 1.38,
+ 1.44, 1.5, 1.56, 1.62, 1.68, 1.74,
+ 1.8, 1.86, 1.92, 1.98, 2.04, 2.1,
+ 2.16, 2.22, 2.28, 2.34, 2.4, 2.46,
+ 2.52, 2.58, 2.64, 2.7, 2.76, 2.82,
+ 2.88, 2.94, 3, 3.06, 3.12, 3.18,
+ 3.24, 3.3, 3.36, 3.42, 3.48, 3.54,
+ 3.6)"
+          idata_min="(-2.394, -2.235, -2.075, -1.915, -1.756, -1.596,
+ -1.437, -1.277, -1.118, -0.9586, -0.7993, -0.6403,
+ -0.4841, -0.3375, -0.2096, -0.1333, -0.1135, -0.1032,
+ -0.09427, -0.08574, -0.07761, -0.06996, -0.06286, -0.05631,
+ -0.05017, -0.04422, -0.03837, -0.03258, -0.02687, -0.02127,
+ -0.01578, -0.01053, -0.005574, -0.0009032, 0.003482, 0.007583,
+ 0.0114, 0.01494, 0.0182, 0.02119, 0.0239, 0.02632,
+ 0.02844, 0.03027, 0.03189, 0.03338, 0.03481, 0.0362,
+ 0.03759, 0.03898, 0.04039, 0.04181, 0.04324, 0.0447,
+ 0.04617, 0.04766, 0.04918, 0.05073, 0.0523, 0.0539,
+ 0.05554, 0.05721, 0.05887, 0.06051, 0.06215, 0.06379,
+ 0.06553, 0.06774, 0.07132, 0.07727, 0.08581, 0.09653,
+ 0.109, 0.1233, 0.143, 0.1988, 0.4466, 0.8356,
+ 1.244, 1.664, 2.088, 2.513, 2.938, 3.364,
+ 3.79, 4.216, 4.641, 5.067, 5.493, 5.919,
+ 6.346)"
+          tdata_0to1_max="(7.19709e-011, 7.82209e-011, 8.44709e-011, 9.07209e-011, 9.69709e-011, 1.03221e-010,
+ 1.09471e-010, 1.15721e-010, 1.21971e-010, 1.28221e-010, 1.34471e-010, 1.40721e-010,
+ 1.46971e-010, 1.53221e-010, 1.59471e-010, 1.65721e-010, 1.71971e-010, 1.78221e-010,
+ 1.84471e-010, 1.90721e-010, 1.96971e-010, 2.03221e-010, 2.09471e-010, 2.15721e-010,
+ 2.21971e-010, 2.28221e-010, 2.34471e-010, 2.40721e-010, 2.46971e-010, 2.53221e-010,
+ 2.59471e-010, 2.65721e-010, 2.71971e-010, 2.78221e-010, 2.84471e-010, 2.90721e-010,
+ 2.96971e-010, 3.03221e-010, 3.09471e-010, 3.15721e-010, 3.21971e-010, 3.28221e-010,
+ 3.34471e-010, 3.40721e-010, 3.46971e-010, 3.53221e-010, 3.59471e-010, 3.65721e-010,
+ 3.71971e-010, 3.78221e-010, 3.84471e-010, 3.90721e-010, 3.96971e-010, 4.03221e-010,
+ 4.09471e-010, 4.15721e-010, 4.21971e-010, 4.28221e-010, 4.34471e-010, 4.40721e-010,
+ 4.46971e-010, 4.53221e-010, 4.59471e-010, 4.65721e-010, 4.71971e-010, 4.78221e-010,
+ 4.84471e-010, 4.90721e-010, 4.96971e-010, 5.03221e-010, 5.09471e-010, 5.15721e-010,
+ 5.21971e-010, 5.28221e-010, 5.34471e-010, 5.40721e-010, 5.46971e-010, 5.53221e-010,
+ 5.59471e-010, 5.65721e-010, 5.71971e-010, 5.78221e-010, 5.84471e-010, 5.90721e-010,
+ 5.96971e-010, 6.03221e-010, 6.09471e-010, 6.15721e-010, 6.21971e-010, 6.28221e-010,
+ 6.34471e-010, 6.40721e-010, 6.46971e-010, 6.53221e-010, 6.59471e-010, 6.65721e-010,
+ 6.71971e-010, 6.78221e-010, 6.84471e-010, 6.90721e-010, 6.96971e-010, 7.03221e-010,
+ 7.09471e-010, 7.15721e-010, 7.21971e-010, 7.28221e-010, 7.34471e-010, 7.40721e-010,
+ 7.46971e-010, 7.53221e-010, 7.59471e-010, 7.65721e-010, 7.71971e-010, 7.78221e-010,
+ 7.84471e-010, 7.90721e-010, 7.96971e-010, 8.03221e-010, 8.09471e-010, 8.15721e-010,
+ 8.21971e-010, 8.28221e-010, 8.34471e-010, 8.40721e-010, 8.46971e-010, 8.53221e-010,
+ 8.59471e-010, 8.65721e-010, 8.71971e-010, 8.78221e-010, 8.84471e-010, 8.90721e-010,
+ 8.96971e-010, 9.03221e-010, 9.09471e-010, 9.15721e-010, 9.21971e-010, 9.28221e-010,
+ 9.34471e-010, 9.40721e-010, 9.46971e-010, 9.53221e-010, 9.59471e-010, 9.65721e-010,
+ 9.71971e-010, 9.78221e-010, 9.84471e-010, 9.90721e-010, 9.96971e-010, 1.00322e-009,
+ 1.00947e-009, 1.01572e-009, 1.02197e-009, 1.02822e-009, 1.03447e-009, 1.04072e-009,
+ 1.04697e-009, 1.05322e-009, 1.05947e-009, 1.06572e-009, 1.07197e-009, 1.07822e-009,
+ 1.08447e-009, 1.09072e-009, 1.09697e-009, 1.10322e-009, 1.10947e-009, 1.11572e-009,
+ 1.12197e-009, 1.12822e-009, 1.13447e-009, 1.14072e-009, 1.14697e-009, 1.15322e-009,
+ 1.15947e-009, 1.16572e-009, 1.17197e-009, 1.17822e-009, 1.18447e-009, 1.19072e-009,
+ 1.19697e-009, 1.20322e-009, 1.20947e-009, 1.21572e-009, 1.22197e-009, 1.22822e-009,
+ 1.23447e-009, 1.24072e-009, 1.24697e-009, 1.25322e-009, 1.25947e-009, 1.26572e-009,
+ 1.27197e-009, 1.27822e-009, 1.28447e-009, 1.29072e-009, 1.29697e-009, 1.30322e-009,
+ 1.30947e-009, 1.31572e-009, 1.32197e-009, 1.32822e-009)"
+          kdata_0to1_max="(0, 0.00144844, 0.00161591, 0.00178283, 0.00194921, 0.00211506,
+ 0.0087038, 0.00937234, 0.0100361, 0.0106951, 0.0113493, 0.0221732,
+ 0.0235462, 0.0248913, 0.0262091, 0.027512, 0.0384896, 0.040387,
+ 0.0422566, 0.0440992, 0.0459152, 0.0477052, 0.0909226, 0.0947716,
+ 0.0985008, 0.102115, 0.10562, 0.151672, 0.156561, 0.161263,
+ 0.165788, 0.170143, 0.231451, 0.237879, 0.244041, 0.249991,
+ 0.255738, 0.306646, 0.314487, 0.322133, 0.329544, 0.346723,
+ 0.354268, 0.361647, 0.368849, 0.375871, 0.436727, 0.446473,
+ 0.456075, 0.465528, 0.47489, 0.508024, 0.518296, 0.528421,
+ 0.538431, 0.548284, 0.578952, 0.589365, 0.599555, 0.609511,
+ 0.619187, 0.661993, 0.673295, 0.684356, 0.695153, 0.695174,
+ 0.703634, 0.711667, 0.719248, 0.725866, 0.705895, 0.708557,
+ 0.710598, 0.711564, 0.710588, 0.813801, 0.819259, 0.824199,
+ 0.827163, 0.82912, 0.854347, 0.858385, 0.861996, 0.865003,
+ 0.86646, 0.82184, 0.821897, 0.821674, 0.821592, 0.821429,
+ 0.86842, 0.871631, 0.874676, 0.877554, 0.928498, 0.936229,
+ 0.943903, 0.951517, 0.95907, 0.902802, 0.908617, 0.914903,
+ 0.921194, 0.927466, 0.912617, 0.919099, 0.925592, 0.932094,
+ 0.938605, 0.915914, 0.921739, 0.928803, 0.935927, 0.943095,
+ 0.982139, 0.992066, 1, 1, 0.970056, 0.977633,
+ 0.985279, 0.992996, 1, 0.981505, 0.988024, 0.995008,
+ 1, 1, 0.97652, 0.981778, 0.987072, 0.992403,
+ 0.997772, 0.989569, 0.994141, 0.99874, 1, 1,
+ 0.958503, 0.959695, 0.960888, 0.961952, 0.984313, 0.987439,
+ 0.99058, 0.993734, 0.996902, 0.986424, 0.988754, 0.991091,
+ 0.993435, 0.995786, 0.984205, 0.985709, 0.987216, 0.988726,
+ 0.990238, 0.991754, 0.993272, 0.994792, 0.996316, 0.997843,
+ 0.997771, 0.99948, 1, 1, 0.978729, 0.978557,
+ 0.978385, 0.978213, 0.978042, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 0.984196, 0.983159, 0.982125, 0.981093, 0.980062,
+ 0.991678, 0.991678, 0.991678, 0.991678, 0.991678, 1,
+ 1, 1, 1, 1)"
+          tdata_1to0_max="(1.63161e-011, 2.2246e-011, 2.81759e-011, 3.41058e-011, 4.00356e-011, 4.59655e-011,
+ 5.18954e-011, 5.78253e-011, 6.37551e-011, 6.9685e-011, 7.56149e-011, 8.15448e-011,
+ 8.74746e-011, 9.34045e-011, 9.93344e-011, 1.05264e-010, 1.11194e-010, 1.17124e-010,
+ 1.23054e-010, 1.28984e-010, 1.34914e-010, 1.40843e-010, 1.46773e-010, 1.52703e-010,
+ 1.58633e-010, 1.64563e-010, 1.70493e-010, 1.76423e-010, 1.82353e-010, 1.88282e-010,
+ 1.94212e-010, 2.00142e-010, 2.06072e-010, 2.12002e-010, 2.17932e-010, 2.23862e-010,
+ 2.29792e-010, 2.35721e-010, 2.41651e-010, 2.47581e-010, 2.53511e-010, 2.59441e-010,
+ 2.65371e-010, 2.71301e-010, 2.77231e-010, 2.8316e-010, 2.8909e-010, 2.9502e-010,
+ 3.0095e-010, 3.0688e-010, 3.1281e-010, 3.1874e-010, 3.2467e-010, 3.30599e-010,
+ 3.36529e-010, 3.42459e-010, 3.48389e-010, 3.54319e-010, 3.60249e-010, 3.66179e-010,
+ 3.72109e-010, 3.78038e-010, 3.83968e-010, 3.89898e-010, 3.95828e-010, 4.01758e-010,
+ 4.07688e-010, 4.13618e-010, 4.19548e-010, 4.25477e-010, 4.31407e-010, 4.37337e-010,
+ 4.43267e-010, 4.49197e-010, 4.55127e-010, 4.61057e-010, 4.66987e-010, 4.72916e-010,
+ 4.78846e-010, 4.84776e-010, 4.90706e-010, 4.96636e-010, 5.02566e-010, 5.08496e-010,
+ 5.14426e-010, 5.20355e-010, 5.26285e-010, 5.32215e-010, 5.38145e-010, 5.44075e-010,
+ 5.50005e-010, 5.55935e-010, 5.61865e-010, 5.67794e-010, 5.73724e-010, 5.79654e-010,
+ 5.85584e-010, 5.91514e-010, 5.97444e-010, 6.03374e-010, 6.09304e-010, 6.15233e-010,
+ 6.21163e-010, 6.27093e-010, 6.33023e-010, 6.38953e-010, 6.44883e-010, 6.50813e-010,
+ 6.56743e-010, 6.62672e-010, 6.68602e-010, 6.74532e-010, 6.80462e-010, 6.86392e-010,
+ 6.92322e-010, 6.98252e-010, 7.04182e-010, 7.10111e-010, 7.16041e-010, 7.21971e-010,
+ 7.27901e-010, 7.33831e-010, 7.39761e-010, 7.45691e-010, 7.51621e-010, 7.5755e-010,
+ 7.6348e-010, 7.6941e-010, 7.7534e-010, 7.8127e-010, 7.872e-010, 7.9313e-010,
+ 7.9906e-010, 8.04989e-010, 8.10919e-010, 8.16849e-010, 8.22779e-010, 8.28709e-010,
+ 8.34639e-010, 8.40569e-010, 8.46499e-010, 8.52428e-010, 8.58358e-010, 8.64288e-010,
+ 8.70218e-010, 8.76148e-010, 8.82078e-010, 8.88008e-010, 8.93938e-010, 8.99867e-010,
+ 9.05797e-010, 9.11727e-010, 9.17657e-010, 9.23587e-010, 9.29517e-010, 9.35447e-010,
+ 9.41377e-010, 9.47306e-010, 9.53236e-010, 9.59166e-010, 9.65096e-010, 9.71026e-010,
+ 9.76956e-010, 9.82886e-010, 9.88816e-010, 9.94745e-010, 1.00068e-009, 1.00661e-009,
+ 1.01254e-009, 1.01846e-009, 1.02439e-009, 1.03032e-009, 1.03625e-009, 1.04218e-009,
+ 1.04811e-009, 1.05404e-009, 1.05997e-009, 1.0659e-009, 1.07183e-009, 1.07776e-009,
+ 1.08369e-009, 1.08962e-009, 1.09555e-009, 1.10148e-009, 1.10741e-009, 1.11334e-009,
+ 1.11927e-009, 1.1252e-009, 1.13113e-009, 1.13706e-009, 1.14299e-009, 1.14892e-009,
+ 1.15485e-009, 1.16078e-009, 1.16671e-009, 1.17264e-009, 1.17857e-009, 1.1845e-009,
+ 1.19043e-009, 1.19636e-009, 1.20229e-009, 1.20822e-009)"
+          kdata_1to0_max="(1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 0.944958, 0.941817, 0.939014,
+ 0.936329, 0.933652, 0.928097, 0.926197, 0.924296, 0.922394,
+ 0.920489, 0.918327, 0.916081, 0.742328, 0.734287, 0.726279,
+ 0.718306, 0.710366, 0.5818, 0.572814, 0.563786, 0.554718,
+ 0.545614, 0.432759, 0.422287, 0.411632, 0.400804, 0.390031,
+ 0.357675, 0.345405, 0.33285, 0.319786, 0.306318, 0.299028,
+ 0.281999, 0.263834, 0.245179, 0.224, 0.21373, 0.19043,
+ 0.164822, 0.138767, 0.11283, 0.168453, 0.142421, 0.11653,
+ 0.0898447, 0.064093, 0.12499, 0.101151, 0.0779349, 0.0556811,
+ 0.0329568, 0.116942, 0.0977118, 0.0785584, 0.0587776, 0.0393621,
+ 0.100619, 0.0856291, 0.0698708, 0.0543328, 0.0388455, 0.0738995,
+ 0.0617298, 0.0492707, 0.0366203, 0.0238299, 0.0109021, 0.0561065,
+ 0.0467763, 0.0372812, 0.0274446, 0.0172799, 0.0457196, 0.0381295,
+ 0.0304268, 0.0225745, 0.0145697, 0.0383468, 0.0325389, 0.0266255,
+ 0.0206042, 0.0144643, 0.0365308, 0.0322321, 0.0277894, 0.0232542,
+ 0.0186239, 0.028672, 0.025203, 0.0216809, 0.0181047, 0.0144733,
+ 0.0148853, 0.0116153, 0.00831567, 0.00498609, 0.0016262, 0.0188761,
+ 0.0170186, 0.015139, 0.0132368, 0.0113117, 0.0155086, 0.0140556,
+ 0.0125899, 0.0111111, 0.00961925, 0.0139533, 0.0129102, 0.0118597,
+ 0.0108016, 0.00973602, 0.0114324, 0.0105801, 0.00972376, 0.00886338,
+ 0.00799891, 0.00901914, 0.00830074, 0.00758063, 0.0068588, 0.00613525,
+ 0.00561266, 0.00490209, 0.00419006, 0.00347656, 0.00276158, 0.00173159,
+ 0.000988725, 0.000244458, 0, 0, 0.00391781, 0.00364127,
+ 0.00336415, 0.00308644, 0.00280814, 0.00360153, 0.003408, 0.00321424,
+ 0.00302027, 0.00282607, 0.00282379, 0.00264561, 0.00246717, 0.00228846,
+ 0.00210949, 0.00204093, 0.00187022, 0.00169929, 0.00152814, 0.00135675,
+ 0.00118514, 0.00121595, 0.00106019, 0.000904174, 0.000747895, 0.000591352,
+ 0.00127719, 0.00118284, 0.00108844, 0.000993996, 0.000899505, 0.000727513,
+ 0.000625664, 0.000523821, 0.000421982, 0.000320148, 0.000293503, 0.000198808,
+ 0.000104067, 9.27975e-006, 0, 0.0004531, 0.000407536, 0.000361956,
+ 0.000316359, 0.000270744, 0.000225112, 0)"
+          vdata_max="(-1.8, -1.74, -1.68, -1.62, -1.56, -1.5,
+ -1.44, -1.38, -1.32, -1.26, -1.2, -1.14,
+ -1.08, -1.02, -0.96, -0.9, -0.84, -0.78,
+ -0.72, -0.66, -0.6, -0.54, -0.48, -0.42,
+ -0.36, -0.3, -0.24, -0.18, -0.12, -0.06,
+ 0, 0.06, 0.12, 0.18, 0.24, 0.3,
+ 0.36, 0.42, 0.48, 0.54, 0.6, 0.66,
+ 0.72, 0.78, 0.84, 0.9, 0.96, 1.02,
+ 1.08, 1.14, 1.2, 1.26, 1.32, 1.38,
+ 1.44, 1.5, 1.56, 1.62, 1.68, 1.74,
+ 1.8, 1.86, 1.92, 1.98, 2.04, 2.1,
+ 2.16, 2.22, 2.28, 2.34, 2.4, 2.46,
+ 2.52, 2.58, 2.64, 2.7, 2.76, 2.82,
+ 2.88, 2.94, 3, 3.06, 3.12, 3.18,
+ 3.24, 3.3, 3.36, 3.42, 3.48, 3.54,
+ 3.6)"
+          idata_max="(-2.394, -2.235, -2.075, -1.915, -1.756, -1.596,
+ -1.437, -1.277, -1.118, -0.9586, -0.7993, -0.6403,
+ -0.4841, -0.3375, -0.2096, -0.1333, -0.1135, -0.1032,
+ -0.09427, -0.08574, -0.07761, -0.06996, -0.06286, -0.05631,
+ -0.05017, -0.04422, -0.03837, -0.03258, -0.02687, -0.02127,
+ -0.01578, -0.01053, -0.005574, -0.0009032, 0.003482, 0.007583,
+ 0.0114, 0.01494, 0.0182, 0.02119, 0.0239, 0.02632,
+ 0.02844, 0.03027, 0.03189, 0.03338, 0.03481, 0.0362,
+ 0.03759, 0.03898, 0.04039, 0.04181, 0.04324, 0.0447,
+ 0.04617, 0.04766, 0.04918, 0.05073, 0.0523, 0.0539,
+ 0.05554, 0.05721, 0.05887, 0.06051, 0.06215, 0.06379,
+ 0.06553, 0.06774, 0.07132, 0.07727, 0.08581, 0.09653,
+ 0.109, 0.1233, 0.143, 0.1988, 0.4466, 0.8356,
+ 1.244, 1.664, 2.088, 2.513, 2.938, 3.364,
+ 3.79, 4.216, 4.641, 5.067, 5.493, 5.919,
+ 6.346)"
+ PORT: a_signal
+       a_PuRef
+       d_pullup_control

.model ibis_ktiv(icx_behavioral) MACRO LANG=VHDLAMS LIB=icxbase
.ends MODEL_U5_1

*Define subcircuit for MODEL_U3_2_ip
.subckt MODEL_U3_2_ip a_signal a_control 
VPullUpRef a_PURef 0 1.8
VPullDownRef a_PDRef 0 1e-100


Y_a_control ibis_driver_logic(icx_behavioral)
+ GENERIC: corner="ibis_typ"
+          vmeas_values="( 0.5, 0.5, 0.5 )"
+ PORT: a_control
+       a_gnd
+       d_control

.model ibis_driver_logic(icx_behavioral) MACRO LANG=VHDLAMS LIB=icxbase

X_126 a_signal d_control 0 a_PURef a_PDRef MODEL_U3_2

.ends MODEL_U3_2_ip

*Define subcircuit for MODEL_U3_2
.subckt MODEL_U3_2 a_signal d_control a_gnd a_PURef a_PDRef

C_comp a_signal a_gnd 6e-012

VGCRef a_GCRef 0 0
G_gnd_clamp a_signal a_GCRef table v(a_signal, a_GCRef) = 
+ (-3,0) (1,0) (2,0) 
+ (6,0) 

VPCRef a_PCRef 0 1.8
G_power_clamp a_PCRef a_signal table v(a_PCRef, a_signal) = 
+ (-6,0) (-2,0) (-1,0) 
+ (3,0) 

Y_control ibis_control(icx_behavioral)
+ PORT: d_control
+       d_pullup_control
+       d_pulldown_control

.model ibis_control(icx_behavioral) MACRO LANG=VHDLAMS LIB=icxbase


*IBIS Pulldown tables
Y_PullDown ibis_ktiv(icx_behavioral)
+ GENERIC: corner="ibis_typ"
+          tdata_0to1_typ="(1.63161e-011, 2.2246e-011, 2.81759e-011, 3.41058e-011, 4.00356e-011, 4.59655e-011,
+ 5.18954e-011, 5.78253e-011, 6.37551e-011, 6.9685e-011, 7.56149e-011, 8.15448e-011,
+ 8.74746e-011, 9.34045e-011, 9.93344e-011, 1.05264e-010, 1.11194e-010, 1.17124e-010,
+ 1.23054e-010, 1.28984e-010, 1.34914e-010, 1.40843e-010, 1.46773e-010, 1.52703e-010,
+ 1.58633e-010, 1.64563e-010, 1.70493e-010, 1.76423e-010, 1.82353e-010, 1.88282e-010,
+ 1.94212e-010, 2.00142e-010, 2.06072e-010, 2.12002e-010, 2.17932e-010, 2.23862e-010,
+ 2.29792e-010, 2.35721e-010, 2.41651e-010, 2.47581e-010, 2.53511e-010, 2.59441e-010,
+ 2.65371e-010, 2.71301e-010, 2.77231e-010, 2.8316e-010, 2.8909e-010, 2.9502e-010,
+ 3.0095e-010, 3.0688e-010, 3.1281e-010, 3.1874e-010, 3.2467e-010, 3.30599e-010,
+ 3.36529e-010, 3.42459e-010, 3.48389e-010, 3.54319e-010, 3.60249e-010, 3.66179e-010,
+ 3.72109e-010, 3.78038e-010, 3.83968e-010, 3.89898e-010, 3.95828e-010, 4.01758e-010,
+ 4.07688e-010, 4.13618e-010, 4.19548e-010, 4.25477e-010, 4.31407e-010, 4.37337e-010,
+ 4.43267e-010, 4.49197e-010, 4.55127e-010, 4.61057e-010, 4.66987e-010, 4.72916e-010,
+ 4.78846e-010, 4.84776e-010, 4.90706e-010, 4.96636e-010, 5.02566e-010, 5.08496e-010,
+ 5.14426e-010, 5.20355e-010, 5.26285e-010, 5.32215e-010, 5.38145e-010, 5.44075e-010,
+ 5.50005e-010, 5.55935e-010, 5.61865e-010, 5.67794e-010, 5.73724e-010, 5.79654e-010,
+ 5.85584e-010, 5.91514e-010, 5.97444e-010, 6.03374e-010, 6.09304e-010, 6.15233e-010,
+ 6.21163e-010, 6.27093e-010, 6.33023e-010, 6.38953e-010, 6.44883e-010, 6.50813e-010,
+ 6.56743e-010, 6.62672e-010, 6.68602e-010, 6.74532e-010, 6.80462e-010, 6.86392e-010,
+ 6.92322e-010, 6.98252e-010, 7.04182e-010, 7.10111e-010, 7.16041e-010, 7.21971e-010,
+ 7.27901e-010, 7.33831e-010, 7.39761e-010, 7.45691e-010, 7.51621e-010, 7.5755e-010,
+ 7.6348e-010, 7.6941e-010, 7.7534e-010, 7.8127e-010, 7.872e-010, 7.9313e-010,
+ 7.9906e-010, 8.04989e-010, 8.10919e-010, 8.16849e-010, 8.22779e-010, 8.28709e-010,
+ 8.34639e-010, 8.40569e-010, 8.46499e-010, 8.52428e-010, 8.58358e-010, 8.64288e-010,
+ 8.70218e-010, 8.76148e-010, 8.82078e-010, 8.88008e-010, 8.93938e-010, 8.99867e-010,
+ 9.05797e-010, 9.11727e-010, 9.17657e-010, 9.23587e-010, 9.29517e-010, 9.35447e-010,
+ 9.41377e-010, 9.47306e-010, 9.53236e-010, 9.59166e-010, 9.65096e-010, 9.71026e-010,
+ 9.76956e-010, 9.82886e-010, 9.88816e-010, 9.94745e-010, 1.00068e-009, 1.00661e-009,
+ 1.01254e-009, 1.01846e-009, 1.02439e-009, 1.03032e-009, 1.03625e-009, 1.04218e-009,
+ 1.04811e-009, 1.05404e-009, 1.05997e-009, 1.0659e-009, 1.07183e-009, 1.07776e-009,
+ 1.08369e-009, 1.08962e-009, 1.09555e-009, 1.10148e-009, 1.10741e-009, 1.11334e-009,
+ 1.11927e-009, 1.1252e-009, 1.13113e-009, 1.13706e-009, 1.14299e-009, 1.14892e-009,
+ 1.15485e-009, 1.16078e-009, 1.16671e-009, 1.17264e-009, 1.17857e-009, 1.1845e-009,
+ 1.19043e-009, 1.19636e-009, 1.20229e-009, 1.20822e-009)"
+          kdata_0to1_typ="(0, 0.00693597, 0.00734267, 0.00775038, 0.00815913, 0.00858505,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0.0149774, 0.0168403, 0.0186985, 0.0205519,
+ 0.0224006, 0.0240851, 0.0257124, 0.0534193, 0.0575498, 0.0616171,
+ 0.0656214, 0.069563, 0.102944, 0.109289, 0.1155, 0.121575,
+ 0.127512, 0.185885, 0.194014, 0.201885, 0.209487, 0.216904,
+ 0.262763, 0.270595, 0.278029, 0.284935, 0.291331, 0.389536,
+ 0.397239, 0.403807, 0.409531, 0.41272, 0.458302, 0.460574,
+ 0.460332, 0.45866, 0.456168, 0.521521, 0.519402, 0.516554,
+ 0.512182, 0.507981, 0.562714, 0.560143, 0.557616, 0.556013,
+ 0.55331, 0.659015, 0.662791, 0.666581, 0.669294, 0.672524,
+ 0.716442, 0.724711, 0.731962, 0.740509, 0.749691, 0.739752,
+ 0.749267, 0.759439, 0.770012, 0.780565, 0.791097, 0.79587,
+ 0.809271, 0.822809, 0.836161, 0.849325, 0.834494, 0.847778,
+ 0.862015, 0.876457, 0.891109, 0.864523, 0.877546, 0.890758,
+ 0.904235, 0.918949, 0.917735, 0.932302, 0.946993, 0.961955,
+ 0.977195, 0.924242, 0.935102, 0.946108, 0.957264, 0.968572,
+ 0.909004, 0.915836, 0.922722, 0.929662, 0.936656, 0.952113,
+ 0.960445, 0.968871, 0.977393, 0.986011, 0.960073, 0.966314,
+ 0.972606, 0.97895, 0.985348, 0.970999, 0.976042, 0.98112,
+ 0.986232, 0.991379, 0.972387, 0.975803, 0.979234, 0.98268,
+ 0.986141, 0.967094, 0.968918, 0.970746, 0.972578, 0.974414,
+ 0.973267, 0.97489, 0.976515, 0.978144, 0.979776, 0.98008,
+ 0.981606, 0.983135, 0.984771, 0.986428, 0.984285, 0.985785,
+ 0.987287, 0.988793, 0.990302, 0.982654, 0.983469, 0.984284,
+ 0.9851, 0.985918, 0.989565, 0.990614, 0.991664, 0.992715,
+ 0.993768, 0.993327, 0.994265, 0.995205, 0.996146, 0.997089,
+ 0.998032, 1, 1, 1, 1, 1,
+ 0.99667, 0.997028, 0.997387, 0.997745, 0.998104, 0.993811,
+ 0.993821, 0.99383, 0.99384, 0.993849, 0.998489, 0.998848,
+ 0.999207, 0.999566, 0.999926, 0.998882, 0.999149, 0.999417,
+ 0.999684, 0.999951, 1, 1)"
+          tdata_1to0_typ="(7.19709e-011, 7.82209e-011, 8.44709e-011, 9.07209e-011, 9.69709e-011, 1.03221e-010,
+ 1.09471e-010, 1.15721e-010, 1.21971e-010, 1.28221e-010, 1.34471e-010, 1.40721e-010,
+ 1.46971e-010, 1.53221e-010, 1.59471e-010, 1.65721e-010, 1.71971e-010, 1.78221e-010,
+ 1.84471e-010, 1.90721e-010, 1.96971e-010, 2.03221e-010, 2.09471e-010, 2.15721e-010,
+ 2.21971e-010, 2.28221e-010, 2.34471e-010, 2.40721e-010, 2.46971e-010, 2.53221e-010,
+ 2.59471e-010, 2.65721e-010, 2.71971e-010, 2.78221e-010, 2.84471e-010, 2.90721e-010,
+ 2.96971e-010, 3.03221e-010, 3.09471e-010, 3.15721e-010, 3.21971e-010, 3.28221e-010,
+ 3.34471e-010, 3.40721e-010, 3.46971e-010, 3.53221e-010, 3.59471e-010, 3.65721e-010,
+ 3.71971e-010, 3.78221e-010, 3.84471e-010, 3.90721e-010, 3.96971e-010, 4.03221e-010,
+ 4.09471e-010, 4.15721e-010, 4.21971e-010, 4.28221e-010, 4.34471e-010, 4.40721e-010,
+ 4.46971e-010, 4.53221e-010, 4.59471e-010, 4.65721e-010, 4.71971e-010, 4.78221e-010,
+ 4.84471e-010, 4.90721e-010, 4.96971e-010, 5.03221e-010, 5.09471e-010, 5.15721e-010,
+ 5.21971e-010, 5.28221e-010, 5.34471e-010, 5.40721e-010, 5.46971e-010, 5.53221e-010,
+ 5.59471e-010, 5.65721e-010, 5.71971e-010, 5.78221e-010, 5.84471e-010, 5.90721e-010,
+ 5.96971e-010, 6.03221e-010, 6.09471e-010, 6.15721e-010, 6.21971e-010, 6.28221e-010,
+ 6.34471e-010, 6.40721e-010, 6.46971e-010, 6.53221e-010, 6.59471e-010, 6.65721e-010,
+ 6.71971e-010, 6.78221e-010, 6.84471e-010, 6.90721e-010, 6.96971e-010, 7.03221e-010,
+ 7.09471e-010, 7.15721e-010, 7.21971e-010, 7.28221e-010, 7.34471e-010, 7.40721e-010,
+ 7.46971e-010, 7.53221e-010, 7.59471e-010, 7.65721e-010, 7.71971e-010, 7.78221e-010,
+ 7.84471e-010, 7.90721e-010, 7.96971e-010, 8.03221e-010, 8.09471e-010, 8.15721e-010,
+ 8.21971e-010, 8.28221e-010, 8.34471e-010, 8.40721e-010, 8.46971e-010, 8.53221e-010,
+ 8.59471e-010, 8.65721e-010, 8.71971e-010, 8.78221e-010, 8.84471e-010, 8.90721e-010,
+ 8.96971e-010, 9.03221e-010, 9.09471e-010, 9.15721e-010, 9.21971e-010, 9.28221e-010,
+ 9.34471e-010, 9.40721e-010, 9.46971e-010, 9.53221e-010, 9.59471e-010, 9.65721e-010,
+ 9.71971e-010, 9.78221e-010, 9.84471e-010, 9.90721e-010, 9.96971e-010, 1.00322e-009,
+ 1.00947e-009, 1.01572e-009, 1.02197e-009, 1.02822e-009, 1.03447e-009, 1.04072e-009,
+ 1.04697e-009, 1.05322e-009, 1.05947e-009, 1.06572e-009, 1.07197e-009, 1.07822e-009,
+ 1.08447e-009, 1.09072e-009, 1.09697e-009, 1.10322e-009, 1.10947e-009, 1.11572e-009,
+ 1.12197e-009, 1.12822e-009, 1.13447e-009, 1.14072e-009, 1.14697e-009, 1.15322e-009,
+ 1.15947e-009, 1.16572e-009, 1.17197e-009, 1.17822e-009, 1.18447e-009, 1.19072e-009,
+ 1.19697e-009, 1.20322e-009, 1.20947e-009, 1.21572e-009, 1.22197e-009, 1.22822e-009,
+ 1.23447e-009, 1.24072e-009, 1.24697e-009, 1.25322e-009, 1.25947e-009, 1.26572e-009,
+ 1.27197e-009, 1.27822e-009, 1.28447e-009, 1.29072e-009, 1.29697e-009, 1.30322e-009,
+ 1.30947e-009, 1.31572e-009, 1.32197e-009, 1.32822e-009)"
+          kdata_1to0_typ="(1, 0.969945, 0.967761, 0.965584, 0.963414, 0.961251,
+ 0.922663, 0.917876, 0.913122, 0.908402, 0.903714, 0.851047,
+ 0.843315, 0.835827, 0.828581, 0.821414, 0.777789, 0.768792,
+ 0.759918, 0.751166, 0.742532, 0.734016, 0.55307, 0.537138,
+ 0.52166, 0.506619, 0.491996, 0.366398, 0.350055, 0.334232,
+ 0.318906, 0.304052, 0.267484, 0.253148, 0.23932, 0.225815,
+ 0.212624, 0.239538, 0.228337, 0.217242, 0.206183, 0.204381,
+ 0.194033, 0.183877, 0.173777, 0.163736, 0.198952, 0.190664,
+ 0.182312, 0.1739, 0.165717, 0.170127, 0.16219, 0.154145,
+ 0.146131, 0.138011, 0.141711, 0.13341, 0.124857, 0.116071,
+ 0.107027, 0.153405, 0.145329, 0.136956, 0.128286, 0.11476,
+ 0.103503, 0.0919088, 0.0799865, 0.0670827, 0.0281211, 0.0117597,
+ 0, 0, 0, 0.0834382, 0.0701074, 0.0565091,
+ 0.0408893, 0.0245442, 0.0671925, 0.0543346, 0.0413051, 0.0277456,
+ 0.0127862, 0.00102775, 0, 0, 0, 0,
+ 0.0193647, 0.0104846, 0.00154843, 0, 0.0346995, 0.0293831,
+ 0.0239779, 0.0184849, 0.012905, 0.0133686, 0.00943205, 0.00530731,
+ 0.00108283, 0, 0.00937699, 0.00689617, 0.00437921, 0.00182603,
+ 0, 0.00216168, 0.000431909, 0, 0, 0,
+ 0.0182273, 0.0184874, 0.018742, 0.0189907, 0.0137603, 0.0140486,
+ 0.0143348, 0.014619, 0.0149012, 0.012462, 0.0127637, 0.0131749,
+ 0.0137195, 0.0142671, 0.00858316, 0.00888649, 0.00919061, 0.00949552,
+ 0.00980122, 0.00658873, 0.00668349, 0.00677755, 0.00687091, 0.00696356,
+ 0, 0, 0, 0, 0.0026533, 0.00305218,
+ 0.00345251, 0.00385433, 0.00425764, 0.00128215, 0.00147873, 0.0016757,
+ 0.00187306, 0.00207081, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0.00312929, 0.00354451, 0.00396081, 0.00437819, 0, 0,
+ 0, 0, 0, 0.00283054, 0.00324669, 0.00366393,
+ 0.00408225, 0.00450167, 0.00320158, 0.00351594, 0.00383091, 0.00414651,
+ 0.00446272, 0.00477956, 0.0034087, 0.00361956, 0.0038307, 0.00404212,
+ 0.00425382, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0.00147984,
+ 0.00168904, 0.00189851, 0.00210825, 0)"
+          vdata_typ="(-1.8, -1.74, -1.68, -1.62, -1.56, -1.5,
+ -1.44, -1.38, -1.32, -1.26, -1.2, -1.14,
+ -1.08, -1.02, -0.96, -0.9, -0.84, -0.78,
+ -0.72, -0.66, -0.6, -0.54, -0.48, -0.42,
+ -0.36, -0.3, -0.24, -0.18, -0.12, -0.06,
+ 0, 0.06, 0.12, 0.18, 0.24, 0.3,
+ 0.36, 0.42, 0.48, 0.54, 0.6, 0.66,
+ 0.72, 0.78, 0.84, 0.9, 0.96, 1.02,
+ 1.08, 1.14, 1.2, 1.26, 1.32, 1.38,
+ 1.44, 1.5, 1.56, 1.62, 1.68, 1.74,
+ 1.8, 1.86, 1.92, 1.98, 2.04, 2.1,
+ 2.16, 2.22, 2.28, 2.34, 2.4, 2.46,
+ 2.52, 2.58, 2.64, 2.7, 2.76, 2.82,
+ 2.88, 2.94, 3, 3.06, 3.12, 3.18,
+ 3.24, 3.3, 3.36, 3.42, 3.48, 3.54,
+ 3.6)"
+          idata_typ="(-6.345, -5.918, -5.492, -5.066, -4.64, -4.214,
+ -3.788, -3.363, -2.937, -2.511, -2.086, -1.663,
+ -1.243, -0.8341, -0.4448, -0.196, -0.1389, -0.1177,
+ -0.1018, -0.08764, -0.075, -0.06428, -0.05584, -0.04952,
+ -0.04448, -0.0399, -0.03541, -0.03094, -0.02644, -0.02194,
+ -0.01743, -0.01301, -0.008738, -0.004612, -0.0006315, 0.003204,
+ 0.006895, 0.01044, 0.01383, 0.01707, 0.02014, 0.02303,
+ 0.02573, 0.02821, 0.03045, 0.03244, 0.0342, 0.03576,
+ 0.03718, 0.03853, 0.03986, 0.0412, 0.04257, 0.04398,
+ 0.04543, 0.04695, 0.04854, 0.0502, 0.05195, 0.05377,
+ 0.05569, 0.0577, 0.05975, 0.06183, 0.06393, 0.06606,
+ 0.06826, 0.07067, 0.07359, 0.0773, 0.08184, 0.08709,
+ 0.09294, 0.09942, 0.1074, 0.1257, 0.2032, 0.3338,
+ 0.4821, 0.6392, 0.7982, 0.9575, 1.116, 1.276,
+ 1.435, 1.595, 1.754, 1.914, 2.073, 2.233,
+ 2.392)"
+          tdata_0to1_min="(1.63161e-011, 2.2246e-011, 2.81759e-011, 3.41058e-011, 4.00356e-011, 4.59655e-011,
+ 5.18954e-011, 5.78253e-011, 6.37551e-011, 6.9685e-011, 7.56149e-011, 8.15448e-011,
+ 8.74746e-011, 9.34045e-011, 9.93344e-011, 1.05264e-010, 1.11194e-010, 1.17124e-010,
+ 1.23054e-010, 1.28984e-010, 1.34914e-010, 1.40843e-010, 1.46773e-010, 1.52703e-010,
+ 1.58633e-010, 1.64563e-010, 1.70493e-010, 1.76423e-010, 1.82353e-010, 1.88282e-010,
+ 1.94212e-010, 2.00142e-010, 2.06072e-010, 2.12002e-010, 2.17932e-010, 2.23862e-010,
+ 2.29792e-010, 2.35721e-010, 2.41651e-010, 2.47581e-010, 2.53511e-010, 2.59441e-010,
+ 2.65371e-010, 2.71301e-010, 2.77231e-010, 2.8316e-010, 2.8909e-010, 2.9502e-010,
+ 3.0095e-010, 3.0688e-010, 3.1281e-010, 3.1874e-010, 3.2467e-010, 3.30599e-010,
+ 3.36529e-010, 3.42459e-010, 3.48389e-010, 3.54319e-010, 3.60249e-010, 3.66179e-010,
+ 3.72109e-010, 3.78038e-010, 3.83968e-010, 3.89898e-010, 3.95828e-010, 4.01758e-010,
+ 4.07688e-010, 4.13618e-010, 4.19548e-010, 4.25477e-010, 4.31407e-010, 4.37337e-010,
+ 4.43267e-010, 4.49197e-010, 4.55127e-010, 4.61057e-010, 4.66987e-010, 4.72916e-010,
+ 4.78846e-010, 4.84776e-010, 4.90706e-010, 4.96636e-010, 5.02566e-010, 5.08496e-010,
+ 5.14426e-010, 5.20355e-010, 5.26285e-010, 5.32215e-010, 5.38145e-010, 5.44075e-010,
+ 5.50005e-010, 5.55935e-010, 5.61865e-010, 5.67794e-010, 5.73724e-010, 5.79654e-010,
+ 5.85584e-010, 5.91514e-010, 5.97444e-010, 6.03374e-010, 6.09304e-010, 6.15233e-010,
+ 6.21163e-010, 6.27093e-010, 6.33023e-010, 6.38953e-010, 6.44883e-010, 6.50813e-010,
+ 6.56743e-010, 6.62672e-010, 6.68602e-010, 6.74532e-010, 6.80462e-010, 6.86392e-010,
+ 6.92322e-010, 6.98252e-010, 7.04182e-010, 7.10111e-010, 7.16041e-010, 7.21971e-010,
+ 7.27901e-010, 7.33831e-010, 7.39761e-010, 7.45691e-010, 7.51621e-010, 7.5755e-010,
+ 7.6348e-010, 7.6941e-010, 7.7534e-010, 7.8127e-010, 7.872e-010, 7.9313e-010,
+ 7.9906e-010, 8.04989e-010, 8.10919e-010, 8.16849e-010, 8.22779e-010, 8.28709e-010,
+ 8.34639e-010, 8.40569e-010, 8.46499e-010, 8.52428e-010, 8.58358e-010, 8.64288e-010,
+ 8.70218e-010, 8.76148e-010, 8.82078e-010, 8.88008e-010, 8.93938e-010, 8.99867e-010,
+ 9.05797e-010, 9.11727e-010, 9.17657e-010, 9.23587e-010, 9.29517e-010, 9.35447e-010,
+ 9.41377e-010, 9.47306e-010, 9.53236e-010, 9.59166e-010, 9.65096e-010, 9.71026e-010,
+ 9.76956e-010, 9.82886e-010, 9.88816e-010, 9.94745e-010, 1.00068e-009, 1.00661e-009,
+ 1.01254e-009, 1.01846e-009, 1.02439e-009, 1.03032e-009, 1.03625e-009, 1.04218e-009,
+ 1.04811e-009, 1.05404e-009, 1.05997e-009, 1.0659e-009, 1.07183e-009, 1.07776e-009,
+ 1.08369e-009, 1.08962e-009, 1.09555e-009, 1.10148e-009, 1.10741e-009, 1.11334e-009,
+ 1.11927e-009, 1.1252e-009, 1.13113e-009, 1.13706e-009, 1.14299e-009, 1.14892e-009,
+ 1.15485e-009, 1.16078e-009, 1.16671e-009, 1.17264e-009, 1.17857e-009, 1.1845e-009,
+ 1.19043e-009, 1.19636e-009, 1.20229e-009, 1.20822e-009)"
+          kdata_0to1_min="(0, 0.00693597, 0.00734267, 0.00775038, 0.00815913, 0.00858505,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0.0149774, 0.0168403, 0.0186985, 0.0205519,
+ 0.0224006, 0.0240851, 0.0257124, 0.0534193, 0.0575498, 0.0616171,
+ 0.0656214, 0.069563, 0.102944, 0.109289, 0.1155, 0.121575,
+ 0.127512, 0.185885, 0.194014, 0.201885, 0.209487, 0.216904,
+ 0.262763, 0.270595, 0.278029, 0.284935, 0.291331, 0.389536,
+ 0.397239, 0.403807, 0.409531, 0.41272, 0.458302, 0.460574,
+ 0.460332, 0.45866, 0.456168, 0.521521, 0.519402, 0.516554,
+ 0.512182, 0.507981, 0.562714, 0.560143, 0.557616, 0.556013,
+ 0.55331, 0.659015, 0.662791, 0.666581, 0.669294, 0.672524,
+ 0.716442, 0.724711, 0.731962, 0.740509, 0.749691, 0.739752,
+ 0.749267, 0.759439, 0.770012, 0.780565, 0.791097, 0.79587,
+ 0.809271, 0.822809, 0.836161, 0.849325, 0.834494, 0.847778,
+ 0.862015, 0.876457, 0.891109, 0.864523, 0.877546, 0.890758,
+ 0.904235, 0.918949, 0.917735, 0.932302, 0.946993, 0.961955,
+ 0.977195, 0.924242, 0.935102, 0.946108, 0.957264, 0.968572,
+ 0.909004, 0.915836, 0.922722, 0.929662, 0.936656, 0.952113,
+ 0.960445, 0.968871, 0.977393, 0.986011, 0.960073, 0.966314,
+ 0.972606, 0.97895, 0.985348, 0.970999, 0.976042, 0.98112,
+ 0.986232, 0.991379, 0.972387, 0.975803, 0.979234, 0.98268,
+ 0.986141, 0.967094, 0.968918, 0.970746, 0.972578, 0.974414,
+ 0.973267, 0.97489, 0.976515, 0.978144, 0.979776, 0.98008,
+ 0.981606, 0.983135, 0.984771, 0.986428, 0.984285, 0.985785,
+ 0.987287, 0.988793, 0.990302, 0.982654, 0.983469, 0.984284,
+ 0.9851, 0.985918, 0.989565, 0.990614, 0.991664, 0.992715,
+ 0.993768, 0.993327, 0.994265, 0.995205, 0.996146, 0.997089,
+ 0.998032, 1, 1, 1, 1, 1,
+ 0.99667, 0.997028, 0.997387, 0.997745, 0.998104, 0.993811,
+ 0.993821, 0.99383, 0.99384, 0.993849, 0.998489, 0.998848,
+ 0.999207, 0.999566, 0.999926, 0.998882, 0.999149, 0.999417,
+ 0.999684, 0.999951, 1, 1)"
+          tdata_1to0_min="(7.19709e-011, 7.82209e-011, 8.44709e-011, 9.07209e-011, 9.69709e-011, 1.03221e-010,
+ 1.09471e-010, 1.15721e-010, 1.21971e-010, 1.28221e-010, 1.34471e-010, 1.40721e-010,
+ 1.46971e-010, 1.53221e-010, 1.59471e-010, 1.65721e-010, 1.71971e-010, 1.78221e-010,
+ 1.84471e-010, 1.90721e-010, 1.96971e-010, 2.03221e-010, 2.09471e-010, 2.15721e-010,
+ 2.21971e-010, 2.28221e-010, 2.34471e-010, 2.40721e-010, 2.46971e-010, 2.53221e-010,
+ 2.59471e-010, 2.65721e-010, 2.71971e-010, 2.78221e-010, 2.84471e-010, 2.90721e-010,
+ 2.96971e-010, 3.03221e-010, 3.09471e-010, 3.15721e-010, 3.21971e-010, 3.28221e-010,
+ 3.34471e-010, 3.40721e-010, 3.46971e-010, 3.53221e-010, 3.59471e-010, 3.65721e-010,
+ 3.71971e-010, 3.78221e-010, 3.84471e-010, 3.90721e-010, 3.96971e-010, 4.03221e-010,
+ 4.09471e-010, 4.15721e-010, 4.21971e-010, 4.28221e-010, 4.34471e-010, 4.40721e-010,
+ 4.46971e-010, 4.53221e-010, 4.59471e-010, 4.65721e-010, 4.71971e-010, 4.78221e-010,
+ 4.84471e-010, 4.90721e-010, 4.96971e-010, 5.03221e-010, 5.09471e-010, 5.15721e-010,
+ 5.21971e-010, 5.28221e-010, 5.34471e-010, 5.40721e-010, 5.46971e-010, 5.53221e-010,
+ 5.59471e-010, 5.65721e-010, 5.71971e-010, 5.78221e-010, 5.84471e-010, 5.90721e-010,
+ 5.96971e-010, 6.03221e-010, 6.09471e-010, 6.15721e-010, 6.21971e-010, 6.28221e-010,
+ 6.34471e-010, 6.40721e-010, 6.46971e-010, 6.53221e-010, 6.59471e-010, 6.65721e-010,
+ 6.71971e-010, 6.78221e-010, 6.84471e-010, 6.90721e-010, 6.96971e-010, 7.03221e-010,
+ 7.09471e-010, 7.15721e-010, 7.21971e-010, 7.28221e-010, 7.34471e-010, 7.40721e-010,
+ 7.46971e-010, 7.53221e-010, 7.59471e-010, 7.65721e-010, 7.71971e-010, 7.78221e-010,
+ 7.84471e-010, 7.90721e-010, 7.96971e-010, 8.03221e-010, 8.09471e-010, 8.15721e-010,
+ 8.21971e-010, 8.28221e-010, 8.34471e-010, 8.40721e-010, 8.46971e-010, 8.53221e-010,
+ 8.59471e-010, 8.65721e-010, 8.71971e-010, 8.78221e-010, 8.84471e-010, 8.90721e-010,
+ 8.96971e-010, 9.03221e-010, 9.09471e-010, 9.15721e-010, 9.21971e-010, 9.28221e-010,
+ 9.34471e-010, 9.40721e-010, 9.46971e-010, 9.53221e-010, 9.59471e-010, 9.65721e-010,
+ 9.71971e-010, 9.78221e-010, 9.84471e-010, 9.90721e-010, 9.96971e-010, 1.00322e-009,
+ 1.00947e-009, 1.01572e-009, 1.02197e-009, 1.02822e-009, 1.03447e-009, 1.04072e-009,
+ 1.04697e-009, 1.05322e-009, 1.05947e-009, 1.06572e-009, 1.07197e-009, 1.07822e-009,
+ 1.08447e-009, 1.09072e-009, 1.09697e-009, 1.10322e-009, 1.10947e-009, 1.11572e-009,
+ 1.12197e-009, 1.12822e-009, 1.13447e-009, 1.14072e-009, 1.14697e-009, 1.15322e-009,
+ 1.15947e-009, 1.16572e-009, 1.17197e-009, 1.17822e-009, 1.18447e-009, 1.19072e-009,
+ 1.19697e-009, 1.20322e-009, 1.20947e-009, 1.21572e-009, 1.22197e-009, 1.22822e-009,
+ 1.23447e-009, 1.24072e-009, 1.24697e-009, 1.25322e-009, 1.25947e-009, 1.26572e-009,
+ 1.27197e-009, 1.27822e-009, 1.28447e-009, 1.29072e-009, 1.29697e-009, 1.30322e-009,
+ 1.30947e-009, 1.31572e-009, 1.32197e-009, 1.32822e-009)"
+          kdata_1to0_min="(1, 0.969945, 0.967761, 0.965584, 0.963414, 0.961251,
+ 0.922663, 0.917876, 0.913122, 0.908402, 0.903714, 0.851047,
+ 0.843315, 0.835827, 0.828581, 0.821414, 0.777789, 0.768792,
+ 0.759918, 0.751166, 0.742532, 0.734016, 0.55307, 0.537138,
+ 0.52166, 0.506619, 0.491996, 0.366398, 0.350055, 0.334232,
+ 0.318906, 0.304052, 0.267484, 0.253148, 0.23932, 0.225815,
+ 0.212624, 0.239538, 0.228337, 0.217242, 0.206183, 0.204381,
+ 0.194033, 0.183877, 0.173777, 0.163736, 0.198952, 0.190664,
+ 0.182312, 0.1739, 0.165717, 0.170127, 0.16219, 0.154145,
+ 0.146131, 0.138011, 0.141711, 0.13341, 0.124857, 0.116071,
+ 0.107027, 0.153405, 0.145329, 0.136956, 0.128286, 0.11476,
+ 0.103503, 0.0919088, 0.0799865, 0.0670827, 0.0281211, 0.0117597,
+ 0, 0, 0, 0.0834382, 0.0701074, 0.0565091,
+ 0.0408893, 0.0245442, 0.0671925, 0.0543346, 0.0413051, 0.0277456,
+ 0.0127862, 0.00102775, 0, 0, 0, 0,
+ 0.0193647, 0.0104846, 0.00154843, 0, 0.0346995, 0.0293831,
+ 0.0239779, 0.0184849, 0.012905, 0.0133686, 0.00943205, 0.00530731,
+ 0.00108283, 0, 0.00937699, 0.00689617, 0.00437921, 0.00182603,
+ 0, 0.00216168, 0.000431909, 0, 0, 0,
+ 0.0182273, 0.0184874, 0.018742, 0.0189907, 0.0137603, 0.0140486,
+ 0.0143348, 0.014619, 0.0149012, 0.012462, 0.0127637, 0.0131749,
+ 0.0137195, 0.0142671, 0.00858316, 0.00888649, 0.00919061, 0.00949552,
+ 0.00980122, 0.00658873, 0.00668349, 0.00677755, 0.00687091, 0.00696356,
+ 0, 0, 0, 0, 0.0026533, 0.00305218,
+ 0.00345251, 0.00385433, 0.00425764, 0.00128215, 0.00147873, 0.0016757,
+ 0.00187306, 0.00207081, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0.00312929, 0.00354451, 0.00396081, 0.00437819, 0, 0,
+ 0, 0, 0, 0.00283054, 0.00324669, 0.00366393,
+ 0.00408225, 0.00450167, 0.00320158, 0.00351594, 0.00383091, 0.00414651,
+ 0.00446272, 0.00477956, 0.0034087, 0.00361956, 0.0038307, 0.00404212,
+ 0.00425382, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0.00147984,
+ 0.00168904, 0.00189851, 0.00210825, 0)"
+          vdata_min="(-1.8, -1.74, -1.68, -1.62, -1.56, -1.5,
+ -1.44, -1.38, -1.32, -1.26, -1.2, -1.14,
+ -1.08, -1.02, -0.96, -0.9, -0.84, -0.78,
+ -0.72, -0.66, -0.6, -0.54, -0.48, -0.42,
+ -0.36, -0.3, -0.24, -0.18, -0.12, -0.06,
+ 0, 0.06, 0.12, 0.18, 0.24, 0.3,
+ 0.36, 0.42, 0.48, 0.54, 0.6, 0.66,
+ 0.72, 0.78, 0.84, 0.9, 0.96, 1.02,
+ 1.08, 1.14, 1.2, 1.26, 1.32, 1.38,
+ 1.44, 1.5, 1.56, 1.62, 1.68, 1.74,
+ 1.8, 1.86, 1.92, 1.98, 2.04, 2.1,
+ 2.16, 2.22, 2.28, 2.34, 2.4, 2.46,
+ 2.52, 2.58, 2.64, 2.7, 2.76, 2.82,
+ 2.88, 2.94, 3, 3.06, 3.12, 3.18,
+ 3.24, 3.3, 3.36, 3.42, 3.48, 3.54,
+ 3.6)"
+          idata_min="(-6.345, -5.918, -5.492, -5.066, -4.64, -4.214,
+ -3.788, -3.363, -2.937, -2.511, -2.086, -1.663,
+ -1.243, -0.8341, -0.4448, -0.196, -0.1389, -0.1177,
+ -0.1018, -0.08764, -0.075, -0.06428, -0.05584, -0.04952,
+ -0.04448, -0.0399, -0.03541, -0.03094, -0.02644, -0.02194,
+ -0.01743, -0.01301, -0.008738, -0.004612, -0.0006315, 0.003204,
+ 0.006895, 0.01044, 0.01383, 0.01707, 0.02014, 0.02303,
+ 0.02573, 0.02821, 0.03045, 0.03244, 0.0342, 0.03576,
+ 0.03718, 0.03853, 0.03986, 0.0412, 0.04257, 0.04398,
+ 0.04543, 0.04695, 0.04854, 0.0502, 0.05195, 0.05377,
+ 0.05569, 0.0577, 0.05975, 0.06183, 0.06393, 0.06606,
+ 0.06826, 0.07067, 0.07359, 0.0773, 0.08184, 0.08709,
+ 0.09294, 0.09942, 0.1074, 0.1257, 0.2032, 0.3338,
+ 0.4821, 0.6392, 0.7982, 0.9575, 1.116, 1.276,
+ 1.435, 1.595, 1.754, 1.914, 2.073, 2.233,
+ 2.392)"
+          tdata_0to1_max="(1.63161e-011, 2.2246e-011, 2.81759e-011, 3.41058e-011, 4.00356e-011, 4.59655e-011,
+ 5.18954e-011, 5.78253e-011, 6.37551e-011, 6.9685e-011, 7.56149e-011, 8.15448e-011,
+ 8.74746e-011, 9.34045e-011, 9.93344e-011, 1.05264e-010, 1.11194e-010, 1.17124e-010,
+ 1.23054e-010, 1.28984e-010, 1.34914e-010, 1.40843e-010, 1.46773e-010, 1.52703e-010,
+ 1.58633e-010, 1.64563e-010, 1.70493e-010, 1.76423e-010, 1.82353e-010, 1.88282e-010,
+ 1.94212e-010, 2.00142e-010, 2.06072e-010, 2.12002e-010, 2.17932e-010, 2.23862e-010,
+ 2.29792e-010, 2.35721e-010, 2.41651e-010, 2.47581e-010, 2.53511e-010, 2.59441e-010,
+ 2.65371e-010, 2.71301e-010, 2.77231e-010, 2.8316e-010, 2.8909e-010, 2.9502e-010,
+ 3.0095e-010, 3.0688e-010, 3.1281e-010, 3.1874e-010, 3.2467e-010, 3.30599e-010,
+ 3.36529e-010, 3.42459e-010, 3.48389e-010, 3.54319e-010, 3.60249e-010, 3.66179e-010,
+ 3.72109e-010, 3.78038e-010, 3.83968e-010, 3.89898e-010, 3.95828e-010, 4.01758e-010,
+ 4.07688e-010, 4.13618e-010, 4.19548e-010, 4.25477e-010, 4.31407e-010, 4.37337e-010,
+ 4.43267e-010, 4.49197e-010, 4.55127e-010, 4.61057e-010, 4.66987e-010, 4.72916e-010,
+ 4.78846e-010, 4.84776e-010, 4.90706e-010, 4.96636e-010, 5.02566e-010, 5.08496e-010,
+ 5.14426e-010, 5.20355e-010, 5.26285e-010, 5.32215e-010, 5.38145e-010, 5.44075e-010,
+ 5.50005e-010, 5.55935e-010, 5.61865e-010, 5.67794e-010, 5.73724e-010, 5.79654e-010,
+ 5.85584e-010, 5.91514e-010, 5.97444e-010, 6.03374e-010, 6.09304e-010, 6.15233e-010,
+ 6.21163e-010, 6.27093e-010, 6.33023e-010, 6.38953e-010, 6.44883e-010, 6.50813e-010,
+ 6.56743e-010, 6.62672e-010, 6.68602e-010, 6.74532e-010, 6.80462e-010, 6.86392e-010,
+ 6.92322e-010, 6.98252e-010, 7.04182e-010, 7.10111e-010, 7.16041e-010, 7.21971e-010,
+ 7.27901e-010, 7.33831e-010, 7.39761e-010, 7.45691e-010, 7.51621e-010, 7.5755e-010,
+ 7.6348e-010, 7.6941e-010, 7.7534e-010, 7.8127e-010, 7.872e-010, 7.9313e-010,
+ 7.9906e-010, 8.04989e-010, 8.10919e-010, 8.16849e-010, 8.22779e-010, 8.28709e-010,
+ 8.34639e-010, 8.40569e-010, 8.46499e-010, 8.52428e-010, 8.58358e-010, 8.64288e-010,
+ 8.70218e-010, 8.76148e-010, 8.82078e-010, 8.88008e-010, 8.93938e-010, 8.99867e-010,
+ 9.05797e-010, 9.11727e-010, 9.17657e-010, 9.23587e-010, 9.29517e-010, 9.35447e-010,
+ 9.41377e-010, 9.47306e-010, 9.53236e-010, 9.59166e-010, 9.65096e-010, 9.71026e-010,
+ 9.76956e-010, 9.82886e-010, 9.88816e-010, 9.94745e-010, 1.00068e-009, 1.00661e-009,
+ 1.01254e-009, 1.01846e-009, 1.02439e-009, 1.03032e-009, 1.03625e-009, 1.04218e-009,
+ 1.04811e-009, 1.05404e-009, 1.05997e-009, 1.0659e-009, 1.07183e-009, 1.07776e-009,
+ 1.08369e-009, 1.08962e-009, 1.09555e-009, 1.10148e-009, 1.10741e-009, 1.11334e-009,
+ 1.11927e-009, 1.1252e-009, 1.13113e-009, 1.13706e-009, 1.14299e-009, 1.14892e-009,
+ 1.15485e-009, 1.16078e-009, 1.16671e-009, 1.17264e-009, 1.17857e-009, 1.1845e-009,
+ 1.19043e-009, 1.19636e-009, 1.20229e-009, 1.20822e-009)"
+          kdata_0to1_max="(0, 0.00693597, 0.00734267, 0.00775038, 0.00815913, 0.00858505,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0.0149774, 0.0168403, 0.0186985, 0.0205519,
+ 0.0224006, 0.0240851, 0.0257124, 0.0534193, 0.0575498, 0.0616171,
+ 0.0656214, 0.069563, 0.102944, 0.109289, 0.1155, 0.121575,
+ 0.127512, 0.185885, 0.194014, 0.201885, 0.209487, 0.216904,
+ 0.262763, 0.270595, 0.278029, 0.284935, 0.291331, 0.389536,
+ 0.397239, 0.403807, 0.409531, 0.41272, 0.458302, 0.460574,
+ 0.460332, 0.45866, 0.456168, 0.521521, 0.519402, 0.516554,
+ 0.512182, 0.507981, 0.562714, 0.560143, 0.557616, 0.556013,
+ 0.55331, 0.659015, 0.662791, 0.666581, 0.669294, 0.672524,
+ 0.716442, 0.724711, 0.731962, 0.740509, 0.749691, 0.739752,
+ 0.749267, 0.759439, 0.770012, 0.780565, 0.791097, 0.79587,
+ 0.809271, 0.822809, 0.836161, 0.849325, 0.834494, 0.847778,
+ 0.862015, 0.876457, 0.891109, 0.864523, 0.877546, 0.890758,
+ 0.904235, 0.918949, 0.917735, 0.932302, 0.946993, 0.961955,
+ 0.977195, 0.924242, 0.935102, 0.946108, 0.957264, 0.968572,
+ 0.909004, 0.915836, 0.922722, 0.929662, 0.936656, 0.952113,
+ 0.960445, 0.968871, 0.977393, 0.986011, 0.960073, 0.966314,
+ 0.972606, 0.97895, 0.985348, 0.970999, 0.976042, 0.98112,
+ 0.986232, 0.991379, 0.972387, 0.975803, 0.979234, 0.98268,
+ 0.986141, 0.967094, 0.968918, 0.970746, 0.972578, 0.974414,
+ 0.973267, 0.97489, 0.976515, 0.978144, 0.979776, 0.98008,
+ 0.981606, 0.983135, 0.984771, 0.986428, 0.984285, 0.985785,
+ 0.987287, 0.988793, 0.990302, 0.982654, 0.983469, 0.984284,
+ 0.9851, 0.985918, 0.989565, 0.990614, 0.991664, 0.992715,
+ 0.993768, 0.993327, 0.994265, 0.995205, 0.996146, 0.997089,
+ 0.998032, 1, 1, 1, 1, 1,
+ 0.99667, 0.997028, 0.997387, 0.997745, 0.998104, 0.993811,
+ 0.993821, 0.99383, 0.99384, 0.993849, 0.998489, 0.998848,
+ 0.999207, 0.999566, 0.999926, 0.998882, 0.999149, 0.999417,
+ 0.999684, 0.999951, 1, 1)"
+          tdata_1to0_max="(7.19709e-011, 7.82209e-011, 8.44709e-011, 9.07209e-011, 9.69709e-011, 1.03221e-010,
+ 1.09471e-010, 1.15721e-010, 1.21971e-010, 1.28221e-010, 1.34471e-010, 1.40721e-010,
+ 1.46971e-010, 1.53221e-010, 1.59471e-010, 1.65721e-010, 1.71971e-010, 1.78221e-010,
+ 1.84471e-010, 1.90721e-010, 1.96971e-010, 2.03221e-010, 2.09471e-010, 2.15721e-010,
+ 2.21971e-010, 2.28221e-010, 2.34471e-010, 2.40721e-010, 2.46971e-010, 2.53221e-010,
+ 2.59471e-010, 2.65721e-010, 2.71971e-010, 2.78221e-010, 2.84471e-010, 2.90721e-010,
+ 2.96971e-010, 3.03221e-010, 3.09471e-010, 3.15721e-010, 3.21971e-010, 3.28221e-010,
+ 3.34471e-010, 3.40721e-010, 3.46971e-010, 3.53221e-010, 3.59471e-010, 3.65721e-010,
+ 3.71971e-010, 3.78221e-010, 3.84471e-010, 3.90721e-010, 3.96971e-010, 4.03221e-010,
+ 4.09471e-010, 4.15721e-010, 4.21971e-010, 4.28221e-010, 4.34471e-010, 4.40721e-010,
+ 4.46971e-010, 4.53221e-010, 4.59471e-010, 4.65721e-010, 4.71971e-010, 4.78221e-010,
+ 4.84471e-010, 4.90721e-010, 4.96971e-010, 5.03221e-010, 5.09471e-010, 5.15721e-010,
+ 5.21971e-010, 5.28221e-010, 5.34471e-010, 5.40721e-010, 5.46971e-010, 5.53221e-010,
+ 5.59471e-010, 5.65721e-010, 5.71971e-010, 5.78221e-010, 5.84471e-010, 5.90721e-010,
+ 5.96971e-010, 6.03221e-010, 6.09471e-010, 6.15721e-010, 6.21971e-010, 6.28221e-010,
+ 6.34471e-010, 6.40721e-010, 6.46971e-010, 6.53221e-010, 6.59471e-010, 6.65721e-010,
+ 6.71971e-010, 6.78221e-010, 6.84471e-010, 6.90721e-010, 6.96971e-010, 7.03221e-010,
+ 7.09471e-010, 7.15721e-010, 7.21971e-010, 7.28221e-010, 7.34471e-010, 7.40721e-010,
+ 7.46971e-010, 7.53221e-010, 7.59471e-010, 7.65721e-010, 7.71971e-010, 7.78221e-010,
+ 7.84471e-010, 7.90721e-010, 7.96971e-010, 8.03221e-010, 8.09471e-010, 8.15721e-010,
+ 8.21971e-010, 8.28221e-010, 8.34471e-010, 8.40721e-010, 8.46971e-010, 8.53221e-010,
+ 8.59471e-010, 8.65721e-010, 8.71971e-010, 8.78221e-010, 8.84471e-010, 8.90721e-010,
+ 8.96971e-010, 9.03221e-010, 9.09471e-010, 9.15721e-010, 9.21971e-010, 9.28221e-010,
+ 9.34471e-010, 9.40721e-010, 9.46971e-010, 9.53221e-010, 9.59471e-010, 9.65721e-010,
+ 9.71971e-010, 9.78221e-010, 9.84471e-010, 9.90721e-010, 9.96971e-010, 1.00322e-009,
+ 1.00947e-009, 1.01572e-009, 1.02197e-009, 1.02822e-009, 1.03447e-009, 1.04072e-009,
+ 1.04697e-009, 1.05322e-009, 1.05947e-009, 1.06572e-009, 1.07197e-009, 1.07822e-009,
+ 1.08447e-009, 1.09072e-009, 1.09697e-009, 1.10322e-009, 1.10947e-009, 1.11572e-009,
+ 1.12197e-009, 1.12822e-009, 1.13447e-009, 1.14072e-009, 1.14697e-009, 1.15322e-009,
+ 1.15947e-009, 1.16572e-009, 1.17197e-009, 1.17822e-009, 1.18447e-009, 1.19072e-009,
+ 1.19697e-009, 1.20322e-009, 1.20947e-009, 1.21572e-009, 1.22197e-009, 1.22822e-009,
+ 1.23447e-009, 1.24072e-009, 1.24697e-009, 1.25322e-009, 1.25947e-009, 1.26572e-009,
+ 1.27197e-009, 1.27822e-009, 1.28447e-009, 1.29072e-009, 1.29697e-009, 1.30322e-009,
+ 1.30947e-009, 1.31572e-009, 1.32197e-009, 1.32822e-009)"
+          kdata_1to0_max="(1, 0.969945, 0.967761, 0.965584, 0.963414, 0.961251,
+ 0.922663, 0.917876, 0.913122, 0.908402, 0.903714, 0.851047,
+ 0.843315, 0.835827, 0.828581, 0.821414, 0.777789, 0.768792,
+ 0.759918, 0.751166, 0.742532, 0.734016, 0.55307, 0.537138,
+ 0.52166, 0.506619, 0.491996, 0.366398, 0.350055, 0.334232,
+ 0.318906, 0.304052, 0.267484, 0.253148, 0.23932, 0.225815,
+ 0.212624, 0.239538, 0.228337, 0.217242, 0.206183, 0.204381,
+ 0.194033, 0.183877, 0.173777, 0.163736, 0.198952, 0.190664,
+ 0.182312, 0.1739, 0.165717, 0.170127, 0.16219, 0.154145,
+ 0.146131, 0.138011, 0.141711, 0.13341, 0.124857, 0.116071,
+ 0.107027, 0.153405, 0.145329, 0.136956, 0.128286, 0.11476,
+ 0.103503, 0.0919088, 0.0799865, 0.0670827, 0.0281211, 0.0117597,
+ 0, 0, 0, 0.0834382, 0.0701074, 0.0565091,
+ 0.0408893, 0.0245442, 0.0671925, 0.0543346, 0.0413051, 0.0277456,
+ 0.0127862, 0.00102775, 0, 0, 0, 0,
+ 0.0193647, 0.0104846, 0.00154843, 0, 0.0346995, 0.0293831,
+ 0.0239779, 0.0184849, 0.012905, 0.0133686, 0.00943205, 0.00530731,
+ 0.00108283, 0, 0.00937699, 0.00689617, 0.00437921, 0.00182603,
+ 0, 0.00216168, 0.000431909, 0, 0, 0,
+ 0.0182273, 0.0184874, 0.018742, 0.0189907, 0.0137603, 0.0140486,
+ 0.0143348, 0.014619, 0.0149012, 0.012462, 0.0127637, 0.0131749,
+ 0.0137195, 0.0142671, 0.00858316, 0.00888649, 0.00919061, 0.00949552,
+ 0.00980122, 0.00658873, 0.00668349, 0.00677755, 0.00687091, 0.00696356,
+ 0, 0, 0, 0, 0.0026533, 0.00305218,
+ 0.00345251, 0.00385433, 0.00425764, 0.00128215, 0.00147873, 0.0016757,
+ 0.00187306, 0.00207081, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0.00312929, 0.00354451, 0.00396081, 0.00437819, 0, 0,
+ 0, 0, 0, 0.00283054, 0.00324669, 0.00366393,
+ 0.00408225, 0.00450167, 0.00320158, 0.00351594, 0.00383091, 0.00414651,
+ 0.00446272, 0.00477956, 0.0034087, 0.00361956, 0.0038307, 0.00404212,
+ 0.00425382, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0.00147984,
+ 0.00168904, 0.00189851, 0.00210825, 0)"
+          vdata_max="(-1.8, -1.74, -1.68, -1.62, -1.56, -1.5,
+ -1.44, -1.38, -1.32, -1.26, -1.2, -1.14,
+ -1.08, -1.02, -0.96, -0.9, -0.84, -0.78,
+ -0.72, -0.66, -0.6, -0.54, -0.48, -0.42,
+ -0.36, -0.3, -0.24, -0.18, -0.12, -0.06,
+ 0, 0.06, 0.12, 0.18, 0.24, 0.3,
+ 0.36, 0.42, 0.48, 0.54, 0.6, 0.66,
+ 0.72, 0.78, 0.84, 0.9, 0.96, 1.02,
+ 1.08, 1.14, 1.2, 1.26, 1.32, 1.38,
+ 1.44, 1.5, 1.56, 1.62, 1.68, 1.74,
+ 1.8, 1.86, 1.92, 1.98, 2.04, 2.1,
+ 2.16, 2.22, 2.28, 2.34, 2.4, 2.46,
+ 2.52, 2.58, 2.64, 2.7, 2.76, 2.82,
+ 2.88, 2.94, 3, 3.06, 3.12, 3.18,
+ 3.24, 3.3, 3.36, 3.42, 3.48, 3.54,
+ 3.6)"
+          idata_max="(-6.345, -5.918, -5.492, -5.066, -4.64, -4.214,
+ -3.788, -3.363, -2.937, -2.511, -2.086, -1.663,
+ -1.243, -0.8341, -0.4448, -0.196, -0.1389, -0.1177,
+ -0.1018, -0.08764, -0.075, -0.06428, -0.05584, -0.04952,
+ -0.04448, -0.0399, -0.03541, -0.03094, -0.02644, -0.02194,
+ -0.01743, -0.01301, -0.008738, -0.004612, -0.0006315, 0.003204,
+ 0.006895, 0.01044, 0.01383, 0.01707, 0.02014, 0.02303,
+ 0.02573, 0.02821, 0.03045, 0.03244, 0.0342, 0.03576,
+ 0.03718, 0.03853, 0.03986, 0.0412, 0.04257, 0.04398,
+ 0.04543, 0.04695, 0.04854, 0.0502, 0.05195, 0.05377,
+ 0.05569, 0.0577, 0.05975, 0.06183, 0.06393, 0.06606,
+ 0.06826, 0.07067, 0.07359, 0.0773, 0.08184, 0.08709,
+ 0.09294, 0.09942, 0.1074, 0.1257, 0.2032, 0.3338,
+ 0.4821, 0.6392, 0.7982, 0.9575, 1.116, 1.276,
+ 1.435, 1.595, 1.754, 1.914, 2.073, 2.233,
+ 2.392)"
+ PORT: a_PdRef
+       a_signal
+       d_pulldown_control


*IBIS Pullup tables
Y_PullUp ibis_ktiv(icx_behavioral)
+ GENERIC: corner="ibis_typ"
+          tdata_0to1_typ="(7.19709e-011, 7.82209e-011, 8.44709e-011, 9.07209e-011, 9.69709e-011, 1.03221e-010,
+ 1.09471e-010, 1.15721e-010, 1.21971e-010, 1.28221e-010, 1.34471e-010, 1.40721e-010,
+ 1.46971e-010, 1.53221e-010, 1.59471e-010, 1.65721e-010, 1.71971e-010, 1.78221e-010,
+ 1.84471e-010, 1.90721e-010, 1.96971e-010, 2.03221e-010, 2.09471e-010, 2.15721e-010,
+ 2.21971e-010, 2.28221e-010, 2.34471e-010, 2.40721e-010, 2.46971e-010, 2.53221e-010,
+ 2.59471e-010, 2.65721e-010, 2.71971e-010, 2.78221e-010, 2.84471e-010, 2.90721e-010,
+ 2.96971e-010, 3.03221e-010, 3.09471e-010, 3.15721e-010, 3.21971e-010, 3.28221e-010,
+ 3.34471e-010, 3.40721e-010, 3.46971e-010, 3.53221e-010, 3.59471e-010, 3.65721e-010,
+ 3.71971e-010, 3.78221e-010, 3.84471e-010, 3.90721e-010, 3.96971e-010, 4.03221e-010,
+ 4.09471e-010, 4.15721e-010, 4.21971e-010, 4.28221e-010, 4.34471e-010, 4.40721e-010,
+ 4.46971e-010, 4.53221e-010, 4.59471e-010, 4.65721e-010, 4.71971e-010, 4.78221e-010,
+ 4.84471e-010, 4.90721e-010, 4.96971e-010, 5.03221e-010, 5.09471e-010, 5.15721e-010,
+ 5.21971e-010, 5.28221e-010, 5.34471e-010, 5.40721e-010, 5.46971e-010, 5.53221e-010,
+ 5.59471e-010, 5.65721e-010, 5.71971e-010, 5.78221e-010, 5.84471e-010, 5.90721e-010,
+ 5.96971e-010, 6.03221e-010, 6.09471e-010, 6.15721e-010, 6.21971e-010, 6.28221e-010,
+ 6.34471e-010, 6.40721e-010, 6.46971e-010, 6.53221e-010, 6.59471e-010, 6.65721e-010,
+ 6.71971e-010, 6.78221e-010, 6.84471e-010, 6.90721e-010, 6.96971e-010, 7.03221e-010,
+ 7.09471e-010, 7.15721e-010, 7.21971e-010, 7.28221e-010, 7.34471e-010, 7.40721e-010,
+ 7.46971e-010, 7.53221e-010, 7.59471e-010, 7.65721e-010, 7.71971e-010, 7.78221e-010,
+ 7.84471e-010, 7.90721e-010, 7.96971e-010, 8.03221e-010, 8.09471e-010, 8.15721e-010,
+ 8.21971e-010, 8.28221e-010, 8.34471e-010, 8.40721e-010, 8.46971e-010, 8.53221e-010,
+ 8.59471e-010, 8.65721e-010, 8.71971e-010, 8.78221e-010, 8.84471e-010, 8.90721e-010,
+ 8.96971e-010, 9.03221e-010, 9.09471e-010, 9.15721e-010, 9.21971e-010, 9.28221e-010,
+ 9.34471e-010, 9.40721e-010, 9.46971e-010, 9.53221e-010, 9.59471e-010, 9.65721e-010,
+ 9.71971e-010, 9.78221e-010, 9.84471e-010, 9.90721e-010, 9.96971e-010, 1.00322e-009,
+ 1.00947e-009, 1.01572e-009, 1.02197e-009, 1.02822e-009, 1.03447e-009, 1.04072e-009,
+ 1.04697e-009, 1.05322e-009, 1.05947e-009, 1.06572e-009, 1.07197e-009, 1.07822e-009,
+ 1.08447e-009, 1.09072e-009, 1.09697e-009, 1.10322e-009, 1.10947e-009, 1.11572e-009,
+ 1.12197e-009, 1.12822e-009, 1.13447e-009, 1.14072e-009, 1.14697e-009, 1.15322e-009,
+ 1.15947e-009, 1.16572e-009, 1.17197e-009, 1.17822e-009, 1.18447e-009, 1.19072e-009,
+ 1.19697e-009, 1.20322e-009, 1.20947e-009, 1.21572e-009, 1.22197e-009, 1.22822e-009,
+ 1.23447e-009, 1.24072e-009, 1.24697e-009, 1.25322e-009, 1.25947e-009, 1.26572e-009,
+ 1.27197e-009, 1.27822e-009, 1.28447e-009, 1.29072e-009, 1.29697e-009, 1.30322e-009,
+ 1.30947e-009, 1.31572e-009, 1.32197e-009, 1.32822e-009)"
+          kdata_0to1_typ="(0, 0.00144844, 0.00161591, 0.00178283, 0.00194921, 0.00211506,
+ 0.0087038, 0.00937234, 0.0100361, 0.0106951, 0.0113493, 0.0221732,
+ 0.0235462, 0.0248913, 0.0262091, 0.027512, 0.0384896, 0.040387,
+ 0.0422566, 0.0440992, 0.0459152, 0.0477052, 0.0909226, 0.0947716,
+ 0.0985008, 0.102115, 0.10562, 0.151672, 0.156561, 0.161263,
+ 0.165788, 0.170143, 0.231451, 0.237879, 0.244041, 0.249991,
+ 0.255738, 0.306646, 0.314487, 0.322133, 0.329544, 0.346723,
+ 0.354268, 0.361647, 0.368849, 0.375871, 0.436727, 0.446473,
+ 0.456075, 0.465528, 0.47489, 0.508024, 0.518296, 0.528421,
+ 0.538431, 0.548284, 0.578952, 0.589365, 0.599555, 0.609511,
+ 0.619187, 0.661993, 0.673295, 0.684356, 0.695153, 0.695174,
+ 0.703634, 0.711667, 0.719248, 0.725866, 0.705895, 0.708557,
+ 0.710598, 0.711564, 0.710588, 0.813801, 0.819259, 0.824199,
+ 0.827163, 0.82912, 0.854347, 0.858385, 0.861996, 0.865003,
+ 0.86646, 0.82184, 0.821897, 0.821674, 0.821592, 0.821429,
+ 0.86842, 0.871631, 0.874676, 0.877554, 0.928498, 0.936229,
+ 0.943903, 0.951517, 0.95907, 0.902802, 0.908617, 0.914903,
+ 0.921194, 0.927466, 0.912617, 0.919099, 0.925592, 0.932094,
+ 0.938605, 0.915914, 0.921739, 0.928803, 0.935927, 0.943095,
+ 0.982139, 0.992066, 1, 1, 0.970056, 0.977633,
+ 0.985279, 0.992996, 1, 0.981505, 0.988024, 0.995008,
+ 1, 1, 0.97652, 0.981778, 0.987072, 0.992403,
+ 0.997772, 0.989569, 0.994141, 0.99874, 1, 1,
+ 0.958503, 0.959695, 0.960888, 0.961952, 0.984313, 0.987439,
+ 0.99058, 0.993734, 0.996902, 0.986424, 0.988754, 0.991091,
+ 0.993435, 0.995786, 0.984205, 0.985709, 0.987216, 0.988726,
+ 0.990238, 0.991754, 0.993272, 0.994792, 0.996316, 0.997843,
+ 0.997771, 0.99948, 1, 1, 0.978729, 0.978557,
+ 0.978385, 0.978213, 0.978042, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 0.984196, 0.983159, 0.982125, 0.981093, 0.980062,
+ 0.991678, 0.991678, 0.991678, 0.991678, 0.991678, 1,
+ 1, 1, 1, 1)"
+          tdata_1to0_typ="(1.63161e-011, 2.2246e-011, 2.81759e-011, 3.41058e-011, 4.00356e-011, 4.59655e-011,
+ 5.18954e-011, 5.78253e-011, 6.37551e-011, 6.9685e-011, 7.56149e-011, 8.15448e-011,
+ 8.74746e-011, 9.34045e-011, 9.93344e-011, 1.05264e-010, 1.11194e-010, 1.17124e-010,
+ 1.23054e-010, 1.28984e-010, 1.34914e-010, 1.40843e-010, 1.46773e-010, 1.52703e-010,
+ 1.58633e-010, 1.64563e-010, 1.70493e-010, 1.76423e-010, 1.82353e-010, 1.88282e-010,
+ 1.94212e-010, 2.00142e-010, 2.06072e-010, 2.12002e-010, 2.17932e-010, 2.23862e-010,
+ 2.29792e-010, 2.35721e-010, 2.41651e-010, 2.47581e-010, 2.53511e-010, 2.59441e-010,
+ 2.65371e-010, 2.71301e-010, 2.77231e-010, 2.8316e-010, 2.8909e-010, 2.9502e-010,
+ 3.0095e-010, 3.0688e-010, 3.1281e-010, 3.1874e-010, 3.2467e-010, 3.30599e-010,
+ 3.36529e-010, 3.42459e-010, 3.48389e-010, 3.54319e-010, 3.60249e-010, 3.66179e-010,
+ 3.72109e-010, 3.78038e-010, 3.83968e-010, 3.89898e-010, 3.95828e-010, 4.01758e-010,
+ 4.07688e-010, 4.13618e-010, 4.19548e-010, 4.25477e-010, 4.31407e-010, 4.37337e-010,
+ 4.43267e-010, 4.49197e-010, 4.55127e-010, 4.61057e-010, 4.66987e-010, 4.72916e-010,
+ 4.78846e-010, 4.84776e-010, 4.90706e-010, 4.96636e-010, 5.02566e-010, 5.08496e-010,
+ 5.14426e-010, 5.20355e-010, 5.26285e-010, 5.32215e-010, 5.38145e-010, 5.44075e-010,
+ 5.50005e-010, 5.55935e-010, 5.61865e-010, 5.67794e-010, 5.73724e-010, 5.79654e-010,
+ 5.85584e-010, 5.91514e-010, 5.97444e-010, 6.03374e-010, 6.09304e-010, 6.15233e-010,
+ 6.21163e-010, 6.27093e-010, 6.33023e-010, 6.38953e-010, 6.44883e-010, 6.50813e-010,
+ 6.56743e-010, 6.62672e-010, 6.68602e-010, 6.74532e-010, 6.80462e-010, 6.86392e-010,
+ 6.92322e-010, 6.98252e-010, 7.04182e-010, 7.10111e-010, 7.16041e-010, 7.21971e-010,
+ 7.27901e-010, 7.33831e-010, 7.39761e-010, 7.45691e-010, 7.51621e-010, 7.5755e-010,
+ 7.6348e-010, 7.6941e-010, 7.7534e-010, 7.8127e-010, 7.872e-010, 7.9313e-010,
+ 7.9906e-010, 8.04989e-010, 8.10919e-010, 8.16849e-010, 8.22779e-010, 8.28709e-010,
+ 8.34639e-010, 8.40569e-010, 8.46499e-010, 8.52428e-010, 8.58358e-010, 8.64288e-010,
+ 8.70218e-010, 8.76148e-010, 8.82078e-010, 8.88008e-010, 8.93938e-010, 8.99867e-010,
+ 9.05797e-010, 9.11727e-010, 9.17657e-010, 9.23587e-010, 9.29517e-010, 9.35447e-010,
+ 9.41377e-010, 9.47306e-010, 9.53236e-010, 9.59166e-010, 9.65096e-010, 9.71026e-010,
+ 9.76956e-010, 9.82886e-010, 9.88816e-010, 9.94745e-010, 1.00068e-009, 1.00661e-009,
+ 1.01254e-009, 1.01846e-009, 1.02439e-009, 1.03032e-009, 1.03625e-009, 1.04218e-009,
+ 1.04811e-009, 1.05404e-009, 1.05997e-009, 1.0659e-009, 1.07183e-009, 1.07776e-009,
+ 1.08369e-009, 1.08962e-009, 1.09555e-009, 1.10148e-009, 1.10741e-009, 1.11334e-009,
+ 1.11927e-009, 1.1252e-009, 1.13113e-009, 1.13706e-009, 1.14299e-009, 1.14892e-009,
+ 1.15485e-009, 1.16078e-009, 1.16671e-009, 1.17264e-009, 1.17857e-009, 1.1845e-009,
+ 1.19043e-009, 1.19636e-009, 1.20229e-009, 1.20822e-009)"
+          kdata_1to0_typ="(1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 0.944958, 0.941817, 0.939014,
+ 0.936329, 0.933652, 0.928097, 0.926197, 0.924296, 0.922394,
+ 0.920489, 0.918327, 0.916081, 0.742328, 0.734287, 0.726279,
+ 0.718306, 0.710366, 0.5818, 0.572814, 0.563786, 0.554718,
+ 0.545614, 0.432759, 0.422287, 0.411632, 0.400804, 0.390031,
+ 0.357675, 0.345405, 0.33285, 0.319786, 0.306318, 0.299028,
+ 0.281999, 0.263834, 0.245179, 0.224, 0.21373, 0.19043,
+ 0.164822, 0.138767, 0.11283, 0.168453, 0.142421, 0.11653,
+ 0.0898447, 0.064093, 0.12499, 0.101151, 0.0779349, 0.0556811,
+ 0.0329568, 0.116942, 0.0977118, 0.0785584, 0.0587776, 0.0393621,
+ 0.100619, 0.0856291, 0.0698708, 0.0543328, 0.0388455, 0.0738995,
+ 0.0617298, 0.0492707, 0.0366203, 0.0238299, 0.0109021, 0.0561065,
+ 0.0467763, 0.0372812, 0.0274446, 0.0172799, 0.0457196, 0.0381295,
+ 0.0304268, 0.0225745, 0.0145697, 0.0383468, 0.0325389, 0.0266255,
+ 0.0206042, 0.0144643, 0.0365308, 0.0322321, 0.0277894, 0.0232542,
+ 0.0186239, 0.028672, 0.025203, 0.0216809, 0.0181047, 0.0144733,
+ 0.0148853, 0.0116153, 0.00831567, 0.00498609, 0.0016262, 0.0188761,
+ 0.0170186, 0.015139, 0.0132368, 0.0113117, 0.0155086, 0.0140556,
+ 0.0125899, 0.0111111, 0.00961925, 0.0139533, 0.0129102, 0.0118597,
+ 0.0108016, 0.00973602, 0.0114324, 0.0105801, 0.00972376, 0.00886338,
+ 0.00799891, 0.00901914, 0.00830074, 0.00758063, 0.0068588, 0.00613525,
+ 0.00561266, 0.00490209, 0.00419006, 0.00347656, 0.00276158, 0.00173159,
+ 0.000988725, 0.000244458, 0, 0, 0.00391781, 0.00364127,
+ 0.00336415, 0.00308644, 0.00280814, 0.00360153, 0.003408, 0.00321424,
+ 0.00302027, 0.00282607, 0.00282379, 0.00264561, 0.00246717, 0.00228846,
+ 0.00210949, 0.00204093, 0.00187022, 0.00169929, 0.00152814, 0.00135675,
+ 0.00118514, 0.00121595, 0.00106019, 0.000904174, 0.000747895, 0.000591352,
+ 0.00127719, 0.00118284, 0.00108844, 0.000993996, 0.000899505, 0.000727513,
+ 0.000625664, 0.000523821, 0.000421982, 0.000320148, 0.000293503, 0.000198808,
+ 0.000104067, 9.27975e-006, 0, 0.0004531, 0.000407536, 0.000361956,
+ 0.000316359, 0.000270744, 0.000225112, 0)"
+          vdata_typ="(-1.8, -1.74, -1.68, -1.62, -1.56, -1.5,
+ -1.44, -1.38, -1.32, -1.26, -1.2, -1.14,
+ -1.08, -1.02, -0.96, -0.9, -0.84, -0.78,
+ -0.72, -0.66, -0.6, -0.54, -0.48, -0.42,
+ -0.36, -0.3, -0.24, -0.18, -0.12, -0.06,
+ 0, 0.06, 0.12, 0.18, 0.24, 0.3,
+ 0.36, 0.42, 0.48, 0.54, 0.6, 0.66,
+ 0.72, 0.78, 0.84, 0.9, 0.96, 1.02,
+ 1.08, 1.14, 1.2, 1.26, 1.32, 1.38,
+ 1.44, 1.5, 1.56, 1.62, 1.68, 1.74,
+ 1.8, 1.86, 1.92, 1.98, 2.04, 2.1,
+ 2.16, 2.22, 2.28, 2.34, 2.4, 2.46,
+ 2.52, 2.58, 2.64, 2.7, 2.76, 2.82,
+ 2.88, 2.94, 3, 3.06, 3.12, 3.18,
+ 3.24, 3.3, 3.36, 3.42, 3.48, 3.54,
+ 3.6)"
+          idata_typ="(-2.394, -2.235, -2.075, -1.915, -1.756, -1.596,
+ -1.437, -1.277, -1.118, -0.9586, -0.7993, -0.6403,
+ -0.4841, -0.3375, -0.2096, -0.1333, -0.1135, -0.1032,
+ -0.09427, -0.08574, -0.07761, -0.06996, -0.06286, -0.05631,
+ -0.05017, -0.04422, -0.03837, -0.03258, -0.02687, -0.02127,
+ -0.01578, -0.01053, -0.005574, -0.0009032, 0.003482, 0.007583,
+ 0.0114, 0.01494, 0.0182, 0.02119, 0.0239, 0.02632,
+ 0.02844, 0.03027, 0.03189, 0.03338, 0.03481, 0.0362,
+ 0.03759, 0.03898, 0.04039, 0.04181, 0.04324, 0.0447,
+ 0.04617, 0.04766, 0.04918, 0.05073, 0.0523, 0.0539,
+ 0.05554, 0.05721, 0.05887, 0.06051, 0.06215, 0.06379,
+ 0.06553, 0.06774, 0.07132, 0.07727, 0.08581, 0.09653,
+ 0.109, 0.1233, 0.143, 0.1988, 0.4466, 0.8356,
+ 1.244, 1.664, 2.088, 2.513, 2.938, 3.364,
+ 3.79, 4.216, 4.641, 5.067, 5.493, 5.919,
+ 6.346)"
+          tdata_0to1_min="(7.19709e-011, 7.82209e-011, 8.44709e-011, 9.07209e-011, 9.69709e-011, 1.03221e-010,
+ 1.09471e-010, 1.15721e-010, 1.21971e-010, 1.28221e-010, 1.34471e-010, 1.40721e-010,
+ 1.46971e-010, 1.53221e-010, 1.59471e-010, 1.65721e-010, 1.71971e-010, 1.78221e-010,
+ 1.84471e-010, 1.90721e-010, 1.96971e-010, 2.03221e-010, 2.09471e-010, 2.15721e-010,
+ 2.21971e-010, 2.28221e-010, 2.34471e-010, 2.40721e-010, 2.46971e-010, 2.53221e-010,
+ 2.59471e-010, 2.65721e-010, 2.71971e-010, 2.78221e-010, 2.84471e-010, 2.90721e-010,
+ 2.96971e-010, 3.03221e-010, 3.09471e-010, 3.15721e-010, 3.21971e-010, 3.28221e-010,
+ 3.34471e-010, 3.40721e-010, 3.46971e-010, 3.53221e-010, 3.59471e-010, 3.65721e-010,
+ 3.71971e-010, 3.78221e-010, 3.84471e-010, 3.90721e-010, 3.96971e-010, 4.03221e-010,
+ 4.09471e-010, 4.15721e-010, 4.21971e-010, 4.28221e-010, 4.34471e-010, 4.40721e-010,
+ 4.46971e-010, 4.53221e-010, 4.59471e-010, 4.65721e-010, 4.71971e-010, 4.78221e-010,
+ 4.84471e-010, 4.90721e-010, 4.96971e-010, 5.03221e-010, 5.09471e-010, 5.15721e-010,
+ 5.21971e-010, 5.28221e-010, 5.34471e-010, 5.40721e-010, 5.46971e-010, 5.53221e-010,
+ 5.59471e-010, 5.65721e-010, 5.71971e-010, 5.78221e-010, 5.84471e-010, 5.90721e-010,
+ 5.96971e-010, 6.03221e-010, 6.09471e-010, 6.15721e-010, 6.21971e-010, 6.28221e-010,
+ 6.34471e-010, 6.40721e-010, 6.46971e-010, 6.53221e-010, 6.59471e-010, 6.65721e-010,
+ 6.71971e-010, 6.78221e-010, 6.84471e-010, 6.90721e-010, 6.96971e-010, 7.03221e-010,
+ 7.09471e-010, 7.15721e-010, 7.21971e-010, 7.28221e-010, 7.34471e-010, 7.40721e-010,
+ 7.46971e-010, 7.53221e-010, 7.59471e-010, 7.65721e-010, 7.71971e-010, 7.78221e-010,
+ 7.84471e-010, 7.90721e-010, 7.96971e-010, 8.03221e-010, 8.09471e-010, 8.15721e-010,
+ 8.21971e-010, 8.28221e-010, 8.34471e-010, 8.40721e-010, 8.46971e-010, 8.53221e-010,
+ 8.59471e-010, 8.65721e-010, 8.71971e-010, 8.78221e-010, 8.84471e-010, 8.90721e-010,
+ 8.96971e-010, 9.03221e-010, 9.09471e-010, 9.15721e-010, 9.21971e-010, 9.28221e-010,
+ 9.34471e-010, 9.40721e-010, 9.46971e-010, 9.53221e-010, 9.59471e-010, 9.65721e-010,
+ 9.71971e-010, 9.78221e-010, 9.84471e-010, 9.90721e-010, 9.96971e-010, 1.00322e-009,
+ 1.00947e-009, 1.01572e-009, 1.02197e-009, 1.02822e-009, 1.03447e-009, 1.04072e-009,
+ 1.04697e-009, 1.05322e-009, 1.05947e-009, 1.06572e-009, 1.07197e-009, 1.07822e-009,
+ 1.08447e-009, 1.09072e-009, 1.09697e-009, 1.10322e-009, 1.10947e-009, 1.11572e-009,
+ 1.12197e-009, 1.12822e-009, 1.13447e-009, 1.14072e-009, 1.14697e-009, 1.15322e-009,
+ 1.15947e-009, 1.16572e-009, 1.17197e-009, 1.17822e-009, 1.18447e-009, 1.19072e-009,
+ 1.19697e-009, 1.20322e-009, 1.20947e-009, 1.21572e-009, 1.22197e-009, 1.22822e-009,
+ 1.23447e-009, 1.24072e-009, 1.24697e-009, 1.25322e-009, 1.25947e-009, 1.26572e-009,
+ 1.27197e-009, 1.27822e-009, 1.28447e-009, 1.29072e-009, 1.29697e-009, 1.30322e-009,
+ 1.30947e-009, 1.31572e-009, 1.32197e-009, 1.32822e-009)"
+          kdata_0to1_min="(0, 0.00144844, 0.00161591, 0.00178283, 0.00194921, 0.00211506,
+ 0.0087038, 0.00937234, 0.0100361, 0.0106951, 0.0113493, 0.0221732,
+ 0.0235462, 0.0248913, 0.0262091, 0.027512, 0.0384896, 0.040387,
+ 0.0422566, 0.0440992, 0.0459152, 0.0477052, 0.0909226, 0.0947716,
+ 0.0985008, 0.102115, 0.10562, 0.151672, 0.156561, 0.161263,
+ 0.165788, 0.170143, 0.231451, 0.237879, 0.244041, 0.249991,
+ 0.255738, 0.306646, 0.314487, 0.322133, 0.329544, 0.346723,
+ 0.354268, 0.361647, 0.368849, 0.375871, 0.436727, 0.446473,
+ 0.456075, 0.465528, 0.47489, 0.508024, 0.518296, 0.528421,
+ 0.538431, 0.548284, 0.578952, 0.589365, 0.599555, 0.609511,
+ 0.619187, 0.661993, 0.673295, 0.684356, 0.695153, 0.695174,
+ 0.703634, 0.711667, 0.719248, 0.725866, 0.705895, 0.708557,
+ 0.710598, 0.711564, 0.710588, 0.813801, 0.819259, 0.824199,
+ 0.827163, 0.82912, 0.854347, 0.858385, 0.861996, 0.865003,
+ 0.86646, 0.82184, 0.821897, 0.821674, 0.821592, 0.821429,
+ 0.86842, 0.871631, 0.874676, 0.877554, 0.928498, 0.936229,
+ 0.943903, 0.951517, 0.95907, 0.902802, 0.908617, 0.914903,
+ 0.921194, 0.927466, 0.912617, 0.919099, 0.925592, 0.932094,
+ 0.938605, 0.915914, 0.921739, 0.928803, 0.935927, 0.943095,
+ 0.982139, 0.992066, 1, 1, 0.970056, 0.977633,
+ 0.985279, 0.992996, 1, 0.981505, 0.988024, 0.995008,
+ 1, 1, 0.97652, 0.981778, 0.987072, 0.992403,
+ 0.997772, 0.989569, 0.994141, 0.99874, 1, 1,
+ 0.958503, 0.959695, 0.960888, 0.961952, 0.984313, 0.987439,
+ 0.99058, 0.993734, 0.996902, 0.986424, 0.988754, 0.991091,
+ 0.993435, 0.995786, 0.984205, 0.985709, 0.987216, 0.988726,
+ 0.990238, 0.991754, 0.993272, 0.994792, 0.996316, 0.997843,
+ 0.997771, 0.99948, 1, 1, 0.978729, 0.978557,
+ 0.978385, 0.978213, 0.978042, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 0.984196, 0.983159, 0.982125, 0.981093, 0.980062,
+ 0.991678, 0.991678, 0.991678, 0.991678, 0.991678, 1,
+ 1, 1, 1, 1)"
+          tdata_1to0_min="(1.63161e-011, 2.2246e-011, 2.81759e-011, 3.41058e-011, 4.00356e-011, 4.59655e-011,
+ 5.18954e-011, 5.78253e-011, 6.37551e-011, 6.9685e-011, 7.56149e-011, 8.15448e-011,
+ 8.74746e-011, 9.34045e-011, 9.93344e-011, 1.05264e-010, 1.11194e-010, 1.17124e-010,
+ 1.23054e-010, 1.28984e-010, 1.34914e-010, 1.40843e-010, 1.46773e-010, 1.52703e-010,
+ 1.58633e-010, 1.64563e-010, 1.70493e-010, 1.76423e-010, 1.82353e-010, 1.88282e-010,
+ 1.94212e-010, 2.00142e-010, 2.06072e-010, 2.12002e-010, 2.17932e-010, 2.23862e-010,
+ 2.29792e-010, 2.35721e-010, 2.41651e-010, 2.47581e-010, 2.53511e-010, 2.59441e-010,
+ 2.65371e-010, 2.71301e-010, 2.77231e-010, 2.8316e-010, 2.8909e-010, 2.9502e-010,
+ 3.0095e-010, 3.0688e-010, 3.1281e-010, 3.1874e-010, 3.2467e-010, 3.30599e-010,
+ 3.36529e-010, 3.42459e-010, 3.48389e-010, 3.54319e-010, 3.60249e-010, 3.66179e-010,
+ 3.72109e-010, 3.78038e-010, 3.83968e-010, 3.89898e-010, 3.95828e-010, 4.01758e-010,
+ 4.07688e-010, 4.13618e-010, 4.19548e-010, 4.25477e-010, 4.31407e-010, 4.37337e-010,
+ 4.43267e-010, 4.49197e-010, 4.55127e-010, 4.61057e-010, 4.66987e-010, 4.72916e-010,
+ 4.78846e-010, 4.84776e-010, 4.90706e-010, 4.96636e-010, 5.02566e-010, 5.08496e-010,
+ 5.14426e-010, 5.20355e-010, 5.26285e-010, 5.32215e-010, 5.38145e-010, 5.44075e-010,
+ 5.50005e-010, 5.55935e-010, 5.61865e-010, 5.67794e-010, 5.73724e-010, 5.79654e-010,
+ 5.85584e-010, 5.91514e-010, 5.97444e-010, 6.03374e-010, 6.09304e-010, 6.15233e-010,
+ 6.21163e-010, 6.27093e-010, 6.33023e-010, 6.38953e-010, 6.44883e-010, 6.50813e-010,
+ 6.56743e-010, 6.62672e-010, 6.68602e-010, 6.74532e-010, 6.80462e-010, 6.86392e-010,
+ 6.92322e-010, 6.98252e-010, 7.04182e-010, 7.10111e-010, 7.16041e-010, 7.21971e-010,
+ 7.27901e-010, 7.33831e-010, 7.39761e-010, 7.45691e-010, 7.51621e-010, 7.5755e-010,
+ 7.6348e-010, 7.6941e-010, 7.7534e-010, 7.8127e-010, 7.872e-010, 7.9313e-010,
+ 7.9906e-010, 8.04989e-010, 8.10919e-010, 8.16849e-010, 8.22779e-010, 8.28709e-010,
+ 8.34639e-010, 8.40569e-010, 8.46499e-010, 8.52428e-010, 8.58358e-010, 8.64288e-010,
+ 8.70218e-010, 8.76148e-010, 8.82078e-010, 8.88008e-010, 8.93938e-010, 8.99867e-010,
+ 9.05797e-010, 9.11727e-010, 9.17657e-010, 9.23587e-010, 9.29517e-010, 9.35447e-010,
+ 9.41377e-010, 9.47306e-010, 9.53236e-010, 9.59166e-010, 9.65096e-010, 9.71026e-010,
+ 9.76956e-010, 9.82886e-010, 9.88816e-010, 9.94745e-010, 1.00068e-009, 1.00661e-009,
+ 1.01254e-009, 1.01846e-009, 1.02439e-009, 1.03032e-009, 1.03625e-009, 1.04218e-009,
+ 1.04811e-009, 1.05404e-009, 1.05997e-009, 1.0659e-009, 1.07183e-009, 1.07776e-009,
+ 1.08369e-009, 1.08962e-009, 1.09555e-009, 1.10148e-009, 1.10741e-009, 1.11334e-009,
+ 1.11927e-009, 1.1252e-009, 1.13113e-009, 1.13706e-009, 1.14299e-009, 1.14892e-009,
+ 1.15485e-009, 1.16078e-009, 1.16671e-009, 1.17264e-009, 1.17857e-009, 1.1845e-009,
+ 1.19043e-009, 1.19636e-009, 1.20229e-009, 1.20822e-009)"
+          kdata_1to0_min="(1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 0.944958, 0.941817, 0.939014,
+ 0.936329, 0.933652, 0.928097, 0.926197, 0.924296, 0.922394,
+ 0.920489, 0.918327, 0.916081, 0.742328, 0.734287, 0.726279,
+ 0.718306, 0.710366, 0.5818, 0.572814, 0.563786, 0.554718,
+ 0.545614, 0.432759, 0.422287, 0.411632, 0.400804, 0.390031,
+ 0.357675, 0.345405, 0.33285, 0.319786, 0.306318, 0.299028,
+ 0.281999, 0.263834, 0.245179, 0.224, 0.21373, 0.19043,
+ 0.164822, 0.138767, 0.11283, 0.168453, 0.142421, 0.11653,
+ 0.0898447, 0.064093, 0.12499, 0.101151, 0.0779349, 0.0556811,
+ 0.0329568, 0.116942, 0.0977118, 0.0785584, 0.0587776, 0.0393621,
+ 0.100619, 0.0856291, 0.0698708, 0.0543328, 0.0388455, 0.0738995,
+ 0.0617298, 0.0492707, 0.0366203, 0.0238299, 0.0109021, 0.0561065,
+ 0.0467763, 0.0372812, 0.0274446, 0.0172799, 0.0457196, 0.0381295,
+ 0.0304268, 0.0225745, 0.0145697, 0.0383468, 0.0325389, 0.0266255,
+ 0.0206042, 0.0144643, 0.0365308, 0.0322321, 0.0277894, 0.0232542,
+ 0.0186239, 0.028672, 0.025203, 0.0216809, 0.0181047, 0.0144733,
+ 0.0148853, 0.0116153, 0.00831567, 0.00498609, 0.0016262, 0.0188761,
+ 0.0170186, 0.015139, 0.0132368, 0.0113117, 0.0155086, 0.0140556,
+ 0.0125899, 0.0111111, 0.00961925, 0.0139533, 0.0129102, 0.0118597,
+ 0.0108016, 0.00973602, 0.0114324, 0.0105801, 0.00972376, 0.00886338,
+ 0.00799891, 0.00901914, 0.00830074, 0.00758063, 0.0068588, 0.00613525,
+ 0.00561266, 0.00490209, 0.00419006, 0.00347656, 0.00276158, 0.00173159,
+ 0.000988725, 0.000244458, 0, 0, 0.00391781, 0.00364127,
+ 0.00336415, 0.00308644, 0.00280814, 0.00360153, 0.003408, 0.00321424,
+ 0.00302027, 0.00282607, 0.00282379, 0.00264561, 0.00246717, 0.00228846,
+ 0.00210949, 0.00204093, 0.00187022, 0.00169929, 0.00152814, 0.00135675,
+ 0.00118514, 0.00121595, 0.00106019, 0.000904174, 0.000747895, 0.000591352,
+ 0.00127719, 0.00118284, 0.00108844, 0.000993996, 0.000899505, 0.000727513,
+ 0.000625664, 0.000523821, 0.000421982, 0.000320148, 0.000293503, 0.000198808,
+ 0.000104067, 9.27975e-006, 0, 0.0004531, 0.000407536, 0.000361956,
+ 0.000316359, 0.000270744, 0.000225112, 0)"
+          vdata_min="(-1.8, -1.74, -1.68, -1.62, -1.56, -1.5,
+ -1.44, -1.38, -1.32, -1.26, -1.2, -1.14,
+ -1.08, -1.02, -0.96, -0.9, -0.84, -0.78,
+ -0.72, -0.66, -0.6, -0.54, -0.48, -0.42,
+ -0.36, -0.3, -0.24, -0.18, -0.12, -0.06,
+ 0, 0.06, 0.12, 0.18, 0.24, 0.3,
+ 0.36, 0.42, 0.48, 0.54, 0.6, 0.66,
+ 0.72, 0.78, 0.84, 0.9, 0.96, 1.02,
+ 1.08, 1.14, 1.2, 1.26, 1.32, 1.38,
+ 1.44, 1.5, 1.56, 1.62, 1.68, 1.74,
+ 1.8, 1.86, 1.92, 1.98, 2.04, 2.1,
+ 2.16, 2.22, 2.28, 2.34, 2.4, 2.46,
+ 2.52, 2.58, 2.64, 2.7, 2.76, 2.82,
+ 2.88, 2.94, 3, 3.06, 3.12, 3.18,
+ 3.24, 3.3, 3.36, 3.42, 3.48, 3.54,
+ 3.6)"
+          idata_min="(-2.394, -2.235, -2.075, -1.915, -1.756, -1.596,
+ -1.437, -1.277, -1.118, -0.9586, -0.7993, -0.6403,
+ -0.4841, -0.3375, -0.2096, -0.1333, -0.1135, -0.1032,
+ -0.09427, -0.08574, -0.07761, -0.06996, -0.06286, -0.05631,
+ -0.05017, -0.04422, -0.03837, -0.03258, -0.02687, -0.02127,
+ -0.01578, -0.01053, -0.005574, -0.0009032, 0.003482, 0.007583,
+ 0.0114, 0.01494, 0.0182, 0.02119, 0.0239, 0.02632,
+ 0.02844, 0.03027, 0.03189, 0.03338, 0.03481, 0.0362,
+ 0.03759, 0.03898, 0.04039, 0.04181, 0.04324, 0.0447,
+ 0.04617, 0.04766, 0.04918, 0.05073, 0.0523, 0.0539,
+ 0.05554, 0.05721, 0.05887, 0.06051, 0.06215, 0.06379,
+ 0.06553, 0.06774, 0.07132, 0.07727, 0.08581, 0.09653,
+ 0.109, 0.1233, 0.143, 0.1988, 0.4466, 0.8356,
+ 1.244, 1.664, 2.088, 2.513, 2.938, 3.364,
+ 3.79, 4.216, 4.641, 5.067, 5.493, 5.919,
+ 6.346)"
+          tdata_0to1_max="(7.19709e-011, 7.82209e-011, 8.44709e-011, 9.07209e-011, 9.69709e-011, 1.03221e-010,
+ 1.09471e-010, 1.15721e-010, 1.21971e-010, 1.28221e-010, 1.34471e-010, 1.40721e-010,
+ 1.46971e-010, 1.53221e-010, 1.59471e-010, 1.65721e-010, 1.71971e-010, 1.78221e-010,
+ 1.84471e-010, 1.90721e-010, 1.96971e-010, 2.03221e-010, 2.09471e-010, 2.15721e-010,
+ 2.21971e-010, 2.28221e-010, 2.34471e-010, 2.40721e-010, 2.46971e-010, 2.53221e-010,
+ 2.59471e-010, 2.65721e-010, 2.71971e-010, 2.78221e-010, 2.84471e-010, 2.90721e-010,
+ 2.96971e-010, 3.03221e-010, 3.09471e-010, 3.15721e-010, 3.21971e-010, 3.28221e-010,
+ 3.34471e-010, 3.40721e-010, 3.46971e-010, 3.53221e-010, 3.59471e-010, 3.65721e-010,
+ 3.71971e-010, 3.78221e-010, 3.84471e-010, 3.90721e-010, 3.96971e-010, 4.03221e-010,
+ 4.09471e-010, 4.15721e-010, 4.21971e-010, 4.28221e-010, 4.34471e-010, 4.40721e-010,
+ 4.46971e-010, 4.53221e-010, 4.59471e-010, 4.65721e-010, 4.71971e-010, 4.78221e-010,
+ 4.84471e-010, 4.90721e-010, 4.96971e-010, 5.03221e-010, 5.09471e-010, 5.15721e-010,
+ 5.21971e-010, 5.28221e-010, 5.34471e-010, 5.40721e-010, 5.46971e-010, 5.53221e-010,
+ 5.59471e-010, 5.65721e-010, 5.71971e-010, 5.78221e-010, 5.84471e-010, 5.90721e-010,
+ 5.96971e-010, 6.03221e-010, 6.09471e-010, 6.15721e-010, 6.21971e-010, 6.28221e-010,
+ 6.34471e-010, 6.40721e-010, 6.46971e-010, 6.53221e-010, 6.59471e-010, 6.65721e-010,
+ 6.71971e-010, 6.78221e-010, 6.84471e-010, 6.90721e-010, 6.96971e-010, 7.03221e-010,
+ 7.09471e-010, 7.15721e-010, 7.21971e-010, 7.28221e-010, 7.34471e-010, 7.40721e-010,
+ 7.46971e-010, 7.53221e-010, 7.59471e-010, 7.65721e-010, 7.71971e-010, 7.78221e-010,
+ 7.84471e-010, 7.90721e-010, 7.96971e-010, 8.03221e-010, 8.09471e-010, 8.15721e-010,
+ 8.21971e-010, 8.28221e-010, 8.34471e-010, 8.40721e-010, 8.46971e-010, 8.53221e-010,
+ 8.59471e-010, 8.65721e-010, 8.71971e-010, 8.78221e-010, 8.84471e-010, 8.90721e-010,
+ 8.96971e-010, 9.03221e-010, 9.09471e-010, 9.15721e-010, 9.21971e-010, 9.28221e-010,
+ 9.34471e-010, 9.40721e-010, 9.46971e-010, 9.53221e-010, 9.59471e-010, 9.65721e-010,
+ 9.71971e-010, 9.78221e-010, 9.84471e-010, 9.90721e-010, 9.96971e-010, 1.00322e-009,
+ 1.00947e-009, 1.01572e-009, 1.02197e-009, 1.02822e-009, 1.03447e-009, 1.04072e-009,
+ 1.04697e-009, 1.05322e-009, 1.05947e-009, 1.06572e-009, 1.07197e-009, 1.07822e-009,
+ 1.08447e-009, 1.09072e-009, 1.09697e-009, 1.10322e-009, 1.10947e-009, 1.11572e-009,
+ 1.12197e-009, 1.12822e-009, 1.13447e-009, 1.14072e-009, 1.14697e-009, 1.15322e-009,
+ 1.15947e-009, 1.16572e-009, 1.17197e-009, 1.17822e-009, 1.18447e-009, 1.19072e-009,
+ 1.19697e-009, 1.20322e-009, 1.20947e-009, 1.21572e-009, 1.22197e-009, 1.22822e-009,
+ 1.23447e-009, 1.24072e-009, 1.24697e-009, 1.25322e-009, 1.25947e-009, 1.26572e-009,
+ 1.27197e-009, 1.27822e-009, 1.28447e-009, 1.29072e-009, 1.29697e-009, 1.30322e-009,
+ 1.30947e-009, 1.31572e-009, 1.32197e-009, 1.32822e-009)"
+          kdata_0to1_max="(0, 0.00144844, 0.00161591, 0.00178283, 0.00194921, 0.00211506,
+ 0.0087038, 0.00937234, 0.0100361, 0.0106951, 0.0113493, 0.0221732,
+ 0.0235462, 0.0248913, 0.0262091, 0.027512, 0.0384896, 0.040387,
+ 0.0422566, 0.0440992, 0.0459152, 0.0477052, 0.0909226, 0.0947716,
+ 0.0985008, 0.102115, 0.10562, 0.151672, 0.156561, 0.161263,
+ 0.165788, 0.170143, 0.231451, 0.237879, 0.244041, 0.249991,
+ 0.255738, 0.306646, 0.314487, 0.322133, 0.329544, 0.346723,
+ 0.354268, 0.361647, 0.368849, 0.375871, 0.436727, 0.446473,
+ 0.456075, 0.465528, 0.47489, 0.508024, 0.518296, 0.528421,
+ 0.538431, 0.548284, 0.578952, 0.589365, 0.599555, 0.609511,
+ 0.619187, 0.661993, 0.673295, 0.684356, 0.695153, 0.695174,
+ 0.703634, 0.711667, 0.719248, 0.725866, 0.705895, 0.708557,
+ 0.710598, 0.711564, 0.710588, 0.813801, 0.819259, 0.824199,
+ 0.827163, 0.82912, 0.854347, 0.858385, 0.861996, 0.865003,
+ 0.86646, 0.82184, 0.821897, 0.821674, 0.821592, 0.821429,
+ 0.86842, 0.871631, 0.874676, 0.877554, 0.928498, 0.936229,
+ 0.943903, 0.951517, 0.95907, 0.902802, 0.908617, 0.914903,
+ 0.921194, 0.927466, 0.912617, 0.919099, 0.925592, 0.932094,
+ 0.938605, 0.915914, 0.921739, 0.928803, 0.935927, 0.943095,
+ 0.982139, 0.992066, 1, 1, 0.970056, 0.977633,
+ 0.985279, 0.992996, 1, 0.981505, 0.988024, 0.995008,
+ 1, 1, 0.97652, 0.981778, 0.987072, 0.992403,
+ 0.997772, 0.989569, 0.994141, 0.99874, 1, 1,
+ 0.958503, 0.959695, 0.960888, 0.961952, 0.984313, 0.987439,
+ 0.99058, 0.993734, 0.996902, 0.986424, 0.988754, 0.991091,
+ 0.993435, 0.995786, 0.984205, 0.985709, 0.987216, 0.988726,
+ 0.990238, 0.991754, 0.993272, 0.994792, 0.996316, 0.997843,
+ 0.997771, 0.99948, 1, 1, 0.978729, 0.978557,
+ 0.978385, 0.978213, 0.978042, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 0.984196, 0.983159, 0.982125, 0.981093, 0.980062,
+ 0.991678, 0.991678, 0.991678, 0.991678, 0.991678, 1,
+ 1, 1, 1, 1)"
+          tdata_1to0_max="(1.63161e-011, 2.2246e-011, 2.81759e-011, 3.41058e-011, 4.00356e-011, 4.59655e-011,
+ 5.18954e-011, 5.78253e-011, 6.37551e-011, 6.9685e-011, 7.56149e-011, 8.15448e-011,
+ 8.74746e-011, 9.34045e-011, 9.93344e-011, 1.05264e-010, 1.11194e-010, 1.17124e-010,
+ 1.23054e-010, 1.28984e-010, 1.34914e-010, 1.40843e-010, 1.46773e-010, 1.52703e-010,
+ 1.58633e-010, 1.64563e-010, 1.70493e-010, 1.76423e-010, 1.82353e-010, 1.88282e-010,
+ 1.94212e-010, 2.00142e-010, 2.06072e-010, 2.12002e-010, 2.17932e-010, 2.23862e-010,
+ 2.29792e-010, 2.35721e-010, 2.41651e-010, 2.47581e-010, 2.53511e-010, 2.59441e-010,
+ 2.65371e-010, 2.71301e-010, 2.77231e-010, 2.8316e-010, 2.8909e-010, 2.9502e-010,
+ 3.0095e-010, 3.0688e-010, 3.1281e-010, 3.1874e-010, 3.2467e-010, 3.30599e-010,
+ 3.36529e-010, 3.42459e-010, 3.48389e-010, 3.54319e-010, 3.60249e-010, 3.66179e-010,
+ 3.72109e-010, 3.78038e-010, 3.83968e-010, 3.89898e-010, 3.95828e-010, 4.01758e-010,
+ 4.07688e-010, 4.13618e-010, 4.19548e-010, 4.25477e-010, 4.31407e-010, 4.37337e-010,
+ 4.43267e-010, 4.49197e-010, 4.55127e-010, 4.61057e-010, 4.66987e-010, 4.72916e-010,
+ 4.78846e-010, 4.84776e-010, 4.90706e-010, 4.96636e-010, 5.02566e-010, 5.08496e-010,
+ 5.14426e-010, 5.20355e-010, 5.26285e-010, 5.32215e-010, 5.38145e-010, 5.44075e-010,
+ 5.50005e-010, 5.55935e-010, 5.61865e-010, 5.67794e-010, 5.73724e-010, 5.79654e-010,
+ 5.85584e-010, 5.91514e-010, 5.97444e-010, 6.03374e-010, 6.09304e-010, 6.15233e-010,
+ 6.21163e-010, 6.27093e-010, 6.33023e-010, 6.38953e-010, 6.44883e-010, 6.50813e-010,
+ 6.56743e-010, 6.62672e-010, 6.68602e-010, 6.74532e-010, 6.80462e-010, 6.86392e-010,
+ 6.92322e-010, 6.98252e-010, 7.04182e-010, 7.10111e-010, 7.16041e-010, 7.21971e-010,
+ 7.27901e-010, 7.33831e-010, 7.39761e-010, 7.45691e-010, 7.51621e-010, 7.5755e-010,
+ 7.6348e-010, 7.6941e-010, 7.7534e-010, 7.8127e-010, 7.872e-010, 7.9313e-010,
+ 7.9906e-010, 8.04989e-010, 8.10919e-010, 8.16849e-010, 8.22779e-010, 8.28709e-010,
+ 8.34639e-010, 8.40569e-010, 8.46499e-010, 8.52428e-010, 8.58358e-010, 8.64288e-010,
+ 8.70218e-010, 8.76148e-010, 8.82078e-010, 8.88008e-010, 8.93938e-010, 8.99867e-010,
+ 9.05797e-010, 9.11727e-010, 9.17657e-010, 9.23587e-010, 9.29517e-010, 9.35447e-010,
+ 9.41377e-010, 9.47306e-010, 9.53236e-010, 9.59166e-010, 9.65096e-010, 9.71026e-010,
+ 9.76956e-010, 9.82886e-010, 9.88816e-010, 9.94745e-010, 1.00068e-009, 1.00661e-009,
+ 1.01254e-009, 1.01846e-009, 1.02439e-009, 1.03032e-009, 1.03625e-009, 1.04218e-009,
+ 1.04811e-009, 1.05404e-009, 1.05997e-009, 1.0659e-009, 1.07183e-009, 1.07776e-009,
+ 1.08369e-009, 1.08962e-009, 1.09555e-009, 1.10148e-009, 1.10741e-009, 1.11334e-009,
+ 1.11927e-009, 1.1252e-009, 1.13113e-009, 1.13706e-009, 1.14299e-009, 1.14892e-009,
+ 1.15485e-009, 1.16078e-009, 1.16671e-009, 1.17264e-009, 1.17857e-009, 1.1845e-009,
+ 1.19043e-009, 1.19636e-009, 1.20229e-009, 1.20822e-009)"
+          kdata_1to0_max="(1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 0.944958, 0.941817, 0.939014,
+ 0.936329, 0.933652, 0.928097, 0.926197, 0.924296, 0.922394,
+ 0.920489, 0.918327, 0.916081, 0.742328, 0.734287, 0.726279,
+ 0.718306, 0.710366, 0.5818, 0.572814, 0.563786, 0.554718,
+ 0.545614, 0.432759, 0.422287, 0.411632, 0.400804, 0.390031,
+ 0.357675, 0.345405, 0.33285, 0.319786, 0.306318, 0.299028,
+ 0.281999, 0.263834, 0.245179, 0.224, 0.21373, 0.19043,
+ 0.164822, 0.138767, 0.11283, 0.168453, 0.142421, 0.11653,
+ 0.0898447, 0.064093, 0.12499, 0.101151, 0.0779349, 0.0556811,
+ 0.0329568, 0.116942, 0.0977118, 0.0785584, 0.0587776, 0.0393621,
+ 0.100619, 0.0856291, 0.0698708, 0.0543328, 0.0388455, 0.0738995,
+ 0.0617298, 0.0492707, 0.0366203, 0.0238299, 0.0109021, 0.0561065,
+ 0.0467763, 0.0372812, 0.0274446, 0.0172799, 0.0457196, 0.0381295,
+ 0.0304268, 0.0225745, 0.0145697, 0.0383468, 0.0325389, 0.0266255,
+ 0.0206042, 0.0144643, 0.0365308, 0.0322321, 0.0277894, 0.0232542,
+ 0.0186239, 0.028672, 0.025203, 0.0216809, 0.0181047, 0.0144733,
+ 0.0148853, 0.0116153, 0.00831567, 0.00498609, 0.0016262, 0.0188761,
+ 0.0170186, 0.015139, 0.0132368, 0.0113117, 0.0155086, 0.0140556,
+ 0.0125899, 0.0111111, 0.00961925, 0.0139533, 0.0129102, 0.0118597,
+ 0.0108016, 0.00973602, 0.0114324, 0.0105801, 0.00972376, 0.00886338,
+ 0.00799891, 0.00901914, 0.00830074, 0.00758063, 0.0068588, 0.00613525,
+ 0.00561266, 0.00490209, 0.00419006, 0.00347656, 0.00276158, 0.00173159,
+ 0.000988725, 0.000244458, 0, 0, 0.00391781, 0.00364127,
+ 0.00336415, 0.00308644, 0.00280814, 0.00360153, 0.003408, 0.00321424,
+ 0.00302027, 0.00282607, 0.00282379, 0.00264561, 0.00246717, 0.00228846,
+ 0.00210949, 0.00204093, 0.00187022, 0.00169929, 0.00152814, 0.00135675,
+ 0.00118514, 0.00121595, 0.00106019, 0.000904174, 0.000747895, 0.000591352,
+ 0.00127719, 0.00118284, 0.00108844, 0.000993996, 0.000899505, 0.000727513,
+ 0.000625664, 0.000523821, 0.000421982, 0.000320148, 0.000293503, 0.000198808,
+ 0.000104067, 9.27975e-006, 0, 0.0004531, 0.000407536, 0.000361956,
+ 0.000316359, 0.000270744, 0.000225112, 0)"
+          vdata_max="(-1.8, -1.74, -1.68, -1.62, -1.56, -1.5,
+ -1.44, -1.38, -1.32, -1.26, -1.2, -1.14,
+ -1.08, -1.02, -0.96, -0.9, -0.84, -0.78,
+ -0.72, -0.66, -0.6, -0.54, -0.48, -0.42,
+ -0.36, -0.3, -0.24, -0.18, -0.12, -0.06,
+ 0, 0.06, 0.12, 0.18, 0.24, 0.3,
+ 0.36, 0.42, 0.48, 0.54, 0.6, 0.66,
+ 0.72, 0.78, 0.84, 0.9, 0.96, 1.02,
+ 1.08, 1.14, 1.2, 1.26, 1.32, 1.38,
+ 1.44, 1.5, 1.56, 1.62, 1.68, 1.74,
+ 1.8, 1.86, 1.92, 1.98, 2.04, 2.1,
+ 2.16, 2.22, 2.28, 2.34, 2.4, 2.46,
+ 2.52, 2.58, 2.64, 2.7, 2.76, 2.82,
+ 2.88, 2.94, 3, 3.06, 3.12, 3.18,
+ 3.24, 3.3, 3.36, 3.42, 3.48, 3.54,
+ 3.6)"
+          idata_max="(-2.394, -2.235, -2.075, -1.915, -1.756, -1.596,
+ -1.437, -1.277, -1.118, -0.9586, -0.7993, -0.6403,
+ -0.4841, -0.3375, -0.2096, -0.1333, -0.1135, -0.1032,
+ -0.09427, -0.08574, -0.07761, -0.06996, -0.06286, -0.05631,
+ -0.05017, -0.04422, -0.03837, -0.03258, -0.02687, -0.02127,
+ -0.01578, -0.01053, -0.005574, -0.0009032, 0.003482, 0.007583,
+ 0.0114, 0.01494, 0.0182, 0.02119, 0.0239, 0.02632,
+ 0.02844, 0.03027, 0.03189, 0.03338, 0.03481, 0.0362,
+ 0.03759, 0.03898, 0.04039, 0.04181, 0.04324, 0.0447,
+ 0.04617, 0.04766, 0.04918, 0.05073, 0.0523, 0.0539,
+ 0.05554, 0.05721, 0.05887, 0.06051, 0.06215, 0.06379,
+ 0.06553, 0.06774, 0.07132, 0.07727, 0.08581, 0.09653,
+ 0.109, 0.1233, 0.143, 0.1988, 0.4466, 0.8356,
+ 1.244, 1.664, 2.088, 2.513, 2.938, 3.364,
+ 3.79, 4.216, 4.641, 5.067, 5.493, 5.919,
+ 6.346)"
+ PORT: a_signal
+       a_PuRef
+       d_pullup_control

.model ibis_ktiv(icx_behavioral) MACRO LANG=VHDLAMS LIB=icxbase
.ends MODEL_U3_2

*Define subcircuit for MODEL_U3_1_ip
.subckt MODEL_U3_1_ip a_signal a_control 
VPullUpRef a_PURef 0 1.8
VPullDownRef a_PDRef 0 1e-100


Y_a_control ibis_driver_logic(icx_behavioral)
+ GENERIC: corner="ibis_typ"
+          vmeas_values="( 0.5, 0.5, 0.5 )"
+ PORT: a_control
+       a_gnd
+       d_control

.model ibis_driver_logic(icx_behavioral) MACRO LANG=VHDLAMS LIB=icxbase

X_136 a_signal d_control 0 a_PURef a_PDRef MODEL_U3_1

.ends MODEL_U3_1_ip

*Define subcircuit for MODEL_U3_1
.subckt MODEL_U3_1 a_signal d_control a_gnd a_PURef a_PDRef

C_comp a_signal a_gnd 6e-012

VGCRef a_GCRef 0 0
G_gnd_clamp a_signal a_GCRef table v(a_signal, a_GCRef) = 
+ (-3,0) (1,0) (2,0) 
+ (6,0) 

VPCRef a_PCRef 0 1.8
G_power_clamp a_PCRef a_signal table v(a_PCRef, a_signal) = 
+ (-6,0) (-2,0) (-1,0) 
+ (3,0) 

Y_control ibis_control(icx_behavioral)
+ PORT: d_control
+       d_pullup_control
+       d_pulldown_control

.model ibis_control(icx_behavioral) MACRO LANG=VHDLAMS LIB=icxbase


*IBIS Pulldown tables
Y_PullDown ibis_ktiv(icx_behavioral)
+ GENERIC: corner="ibis_typ"
+          tdata_0to1_typ="(1.63161e-011, 2.2246e-011, 2.81759e-011, 3.41058e-011, 4.00356e-011, 4.59655e-011,
+ 5.18954e-011, 5.78253e-011, 6.37551e-011, 6.9685e-011, 7.56149e-011, 8.15448e-011,
+ 8.74746e-011, 9.34045e-011, 9.93344e-011, 1.05264e-010, 1.11194e-010, 1.17124e-010,
+ 1.23054e-010, 1.28984e-010, 1.34914e-010, 1.40843e-010, 1.46773e-010, 1.52703e-010,
+ 1.58633e-010, 1.64563e-010, 1.70493e-010, 1.76423e-010, 1.82353e-010, 1.88282e-010,
+ 1.94212e-010, 2.00142e-010, 2.06072e-010, 2.12002e-010, 2.17932e-010, 2.23862e-010,
+ 2.29792e-010, 2.35721e-010, 2.41651e-010, 2.47581e-010, 2.53511e-010, 2.59441e-010,
+ 2.65371e-010, 2.71301e-010, 2.77231e-010, 2.8316e-010, 2.8909e-010, 2.9502e-010,
+ 3.0095e-010, 3.0688e-010, 3.1281e-010, 3.1874e-010, 3.2467e-010, 3.30599e-010,
+ 3.36529e-010, 3.42459e-010, 3.48389e-010, 3.54319e-010, 3.60249e-010, 3.66179e-010,
+ 3.72109e-010, 3.78038e-010, 3.83968e-010, 3.89898e-010, 3.95828e-010, 4.01758e-010,
+ 4.07688e-010, 4.13618e-010, 4.19548e-010, 4.25477e-010, 4.31407e-010, 4.37337e-010,
+ 4.43267e-010, 4.49197e-010, 4.55127e-010, 4.61057e-010, 4.66987e-010, 4.72916e-010,
+ 4.78846e-010, 4.84776e-010, 4.90706e-010, 4.96636e-010, 5.02566e-010, 5.08496e-010,
+ 5.14426e-010, 5.20355e-010, 5.26285e-010, 5.32215e-010, 5.38145e-010, 5.44075e-010,
+ 5.50005e-010, 5.55935e-010, 5.61865e-010, 5.67794e-010, 5.73724e-010, 5.79654e-010,
+ 5.85584e-010, 5.91514e-010, 5.97444e-010, 6.03374e-010, 6.09304e-010, 6.15233e-010,
+ 6.21163e-010, 6.27093e-010, 6.33023e-010, 6.38953e-010, 6.44883e-010, 6.50813e-010,
+ 6.56743e-010, 6.62672e-010, 6.68602e-010, 6.74532e-010, 6.80462e-010, 6.86392e-010,
+ 6.92322e-010, 6.98252e-010, 7.04182e-010, 7.10111e-010, 7.16041e-010, 7.21971e-010,
+ 7.27901e-010, 7.33831e-010, 7.39761e-010, 7.45691e-010, 7.51621e-010, 7.5755e-010,
+ 7.6348e-010, 7.6941e-010, 7.7534e-010, 7.8127e-010, 7.872e-010, 7.9313e-010,
+ 7.9906e-010, 8.04989e-010, 8.10919e-010, 8.16849e-010, 8.22779e-010, 8.28709e-010,
+ 8.34639e-010, 8.40569e-010, 8.46499e-010, 8.52428e-010, 8.58358e-010, 8.64288e-010,
+ 8.70218e-010, 8.76148e-010, 8.82078e-010, 8.88008e-010, 8.93938e-010, 8.99867e-010,
+ 9.05797e-010, 9.11727e-010, 9.17657e-010, 9.23587e-010, 9.29517e-010, 9.35447e-010,
+ 9.41377e-010, 9.47306e-010, 9.53236e-010, 9.59166e-010, 9.65096e-010, 9.71026e-010,
+ 9.76956e-010, 9.82886e-010, 9.88816e-010, 9.94745e-010, 1.00068e-009, 1.00661e-009,
+ 1.01254e-009, 1.01846e-009, 1.02439e-009, 1.03032e-009, 1.03625e-009, 1.04218e-009,
+ 1.04811e-009, 1.05404e-009, 1.05997e-009, 1.0659e-009, 1.07183e-009, 1.07776e-009,
+ 1.08369e-009, 1.08962e-009, 1.09555e-009, 1.10148e-009, 1.10741e-009, 1.11334e-009,
+ 1.11927e-009, 1.1252e-009, 1.13113e-009, 1.13706e-009, 1.14299e-009, 1.14892e-009,
+ 1.15485e-009, 1.16078e-009, 1.16671e-009, 1.17264e-009, 1.17857e-009, 1.1845e-009,
+ 1.19043e-009, 1.19636e-009, 1.20229e-009, 1.20822e-009)"
+          kdata_0to1_typ="(0, 0.00693597, 0.00734267, 0.00775038, 0.00815913, 0.00858505,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0.0149774, 0.0168403, 0.0186985, 0.0205519,
+ 0.0224006, 0.0240851, 0.0257124, 0.0534193, 0.0575498, 0.0616171,
+ 0.0656214, 0.069563, 0.102944, 0.109289, 0.1155, 0.121575,
+ 0.127512, 0.185885, 0.194014, 0.201885, 0.209487, 0.216904,
+ 0.262763, 0.270595, 0.278029, 0.284935, 0.291331, 0.389536,
+ 0.397239, 0.403807, 0.409531, 0.41272, 0.458302, 0.460574,
+ 0.460332, 0.45866, 0.456168, 0.521521, 0.519402, 0.516554,
+ 0.512182, 0.507981, 0.562714, 0.560143, 0.557616, 0.556013,
+ 0.55331, 0.659015, 0.662791, 0.666581, 0.669294, 0.672524,
+ 0.716442, 0.724711, 0.731962, 0.740509, 0.749691, 0.739752,
+ 0.749267, 0.759439, 0.770012, 0.780565, 0.791097, 0.79587,
+ 0.809271, 0.822809, 0.836161, 0.849325, 0.834494, 0.847778,
+ 0.862015, 0.876457, 0.891109, 0.864523, 0.877546, 0.890758,
+ 0.904235, 0.918949, 0.917735, 0.932302, 0.946993, 0.961955,
+ 0.977195, 0.924242, 0.935102, 0.946108, 0.957264, 0.968572,
+ 0.909004, 0.915836, 0.922722, 0.929662, 0.936656, 0.952113,
+ 0.960445, 0.968871, 0.977393, 0.986011, 0.960073, 0.966314,
+ 0.972606, 0.97895, 0.985348, 0.970999, 0.976042, 0.98112,
+ 0.986232, 0.991379, 0.972387, 0.975803, 0.979234, 0.98268,
+ 0.986141, 0.967094, 0.968918, 0.970746, 0.972578, 0.974414,
+ 0.973267, 0.97489, 0.976515, 0.978144, 0.979776, 0.98008,
+ 0.981606, 0.983135, 0.984771, 0.986428, 0.984285, 0.985785,
+ 0.987287, 0.988793, 0.990302, 0.982654, 0.983469, 0.984284,
+ 0.9851, 0.985918, 0.989565, 0.990614, 0.991664, 0.992715,
+ 0.993768, 0.993327, 0.994265, 0.995205, 0.996146, 0.997089,
+ 0.998032, 1, 1, 1, 1, 1,
+ 0.99667, 0.997028, 0.997387, 0.997745, 0.998104, 0.993811,
+ 0.993821, 0.99383, 0.99384, 0.993849, 0.998489, 0.998848,
+ 0.999207, 0.999566, 0.999926, 0.998882, 0.999149, 0.999417,
+ 0.999684, 0.999951, 1, 1)"
+          tdata_1to0_typ="(7.19709e-011, 7.82209e-011, 8.44709e-011, 9.07209e-011, 9.69709e-011, 1.03221e-010,
+ 1.09471e-010, 1.15721e-010, 1.21971e-010, 1.28221e-010, 1.34471e-010, 1.40721e-010,
+ 1.46971e-010, 1.53221e-010, 1.59471e-010, 1.65721e-010, 1.71971e-010, 1.78221e-010,
+ 1.84471e-010, 1.90721e-010, 1.96971e-010, 2.03221e-010, 2.09471e-010, 2.15721e-010,
+ 2.21971e-010, 2.28221e-010, 2.34471e-010, 2.40721e-010, 2.46971e-010, 2.53221e-010,
+ 2.59471e-010, 2.65721e-010, 2.71971e-010, 2.78221e-010, 2.84471e-010, 2.90721e-010,
+ 2.96971e-010, 3.03221e-010, 3.09471e-010, 3.15721e-010, 3.21971e-010, 3.28221e-010,
+ 3.34471e-010, 3.40721e-010, 3.46971e-010, 3.53221e-010, 3.59471e-010, 3.65721e-010,
+ 3.71971e-010, 3.78221e-010, 3.84471e-010, 3.90721e-010, 3.96971e-010, 4.03221e-010,
+ 4.09471e-010, 4.15721e-010, 4.21971e-010, 4.28221e-010, 4.34471e-010, 4.40721e-010,
+ 4.46971e-010, 4.53221e-010, 4.59471e-010, 4.65721e-010, 4.71971e-010, 4.78221e-010,
+ 4.84471e-010, 4.90721e-010, 4.96971e-010, 5.03221e-010, 5.09471e-010, 5.15721e-010,
+ 5.21971e-010, 5.28221e-010, 5.34471e-010, 5.40721e-010, 5.46971e-010, 5.53221e-010,
+ 5.59471e-010, 5.65721e-010, 5.71971e-010, 5.78221e-010, 5.84471e-010, 5.90721e-010,
+ 5.96971e-010, 6.03221e-010, 6.09471e-010, 6.15721e-010, 6.21971e-010, 6.28221e-010,
+ 6.34471e-010, 6.40721e-010, 6.46971e-010, 6.53221e-010, 6.59471e-010, 6.65721e-010,
+ 6.71971e-010, 6.78221e-010, 6.84471e-010, 6.90721e-010, 6.96971e-010, 7.03221e-010,
+ 7.09471e-010, 7.15721e-010, 7.21971e-010, 7.28221e-010, 7.34471e-010, 7.40721e-010,
+ 7.46971e-010, 7.53221e-010, 7.59471e-010, 7.65721e-010, 7.71971e-010, 7.78221e-010,
+ 7.84471e-010, 7.90721e-010, 7.96971e-010, 8.03221e-010, 8.09471e-010, 8.15721e-010,
+ 8.21971e-010, 8.28221e-010, 8.34471e-010, 8.40721e-010, 8.46971e-010, 8.53221e-010,
+ 8.59471e-010, 8.65721e-010, 8.71971e-010, 8.78221e-010, 8.84471e-010, 8.90721e-010,
+ 8.96971e-010, 9.03221e-010, 9.09471e-010, 9.15721e-010, 9.21971e-010, 9.28221e-010,
+ 9.34471e-010, 9.40721e-010, 9.46971e-010, 9.53221e-010, 9.59471e-010, 9.65721e-010,
+ 9.71971e-010, 9.78221e-010, 9.84471e-010, 9.90721e-010, 9.96971e-010, 1.00322e-009,
+ 1.00947e-009, 1.01572e-009, 1.02197e-009, 1.02822e-009, 1.03447e-009, 1.04072e-009,
+ 1.04697e-009, 1.05322e-009, 1.05947e-009, 1.06572e-009, 1.07197e-009, 1.07822e-009,
+ 1.08447e-009, 1.09072e-009, 1.09697e-009, 1.10322e-009, 1.10947e-009, 1.11572e-009,
+ 1.12197e-009, 1.12822e-009, 1.13447e-009, 1.14072e-009, 1.14697e-009, 1.15322e-009,
+ 1.15947e-009, 1.16572e-009, 1.17197e-009, 1.17822e-009, 1.18447e-009, 1.19072e-009,
+ 1.19697e-009, 1.20322e-009, 1.20947e-009, 1.21572e-009, 1.22197e-009, 1.22822e-009,
+ 1.23447e-009, 1.24072e-009, 1.24697e-009, 1.25322e-009, 1.25947e-009, 1.26572e-009,
+ 1.27197e-009, 1.27822e-009, 1.28447e-009, 1.29072e-009, 1.29697e-009, 1.30322e-009,
+ 1.30947e-009, 1.31572e-009, 1.32197e-009, 1.32822e-009)"
+          kdata_1to0_typ="(1, 0.969945, 0.967761, 0.965584, 0.963414, 0.961251,
+ 0.922663, 0.917876, 0.913122, 0.908402, 0.903714, 0.851047,
+ 0.843315, 0.835827, 0.828581, 0.821414, 0.777789, 0.768792,
+ 0.759918, 0.751166, 0.742532, 0.734016, 0.55307, 0.537138,
+ 0.52166, 0.506619, 0.491996, 0.366398, 0.350055, 0.334232,
+ 0.318906, 0.304052, 0.267484, 0.253148, 0.23932, 0.225815,
+ 0.212624, 0.239538, 0.228337, 0.217242, 0.206183, 0.204381,
+ 0.194033, 0.183877, 0.173777, 0.163736, 0.198952, 0.190664,
+ 0.182312, 0.1739, 0.165717, 0.170127, 0.16219, 0.154145,
+ 0.146131, 0.138011, 0.141711, 0.13341, 0.124857, 0.116071,
+ 0.107027, 0.153405, 0.145329, 0.136956, 0.128286, 0.11476,
+ 0.103503, 0.0919088, 0.0799865, 0.0670827, 0.0281211, 0.0117597,
+ 0, 0, 0, 0.0834382, 0.0701074, 0.0565091,
+ 0.0408893, 0.0245442, 0.0671925, 0.0543346, 0.0413051, 0.0277456,
+ 0.0127862, 0.00102775, 0, 0, 0, 0,
+ 0.0193647, 0.0104846, 0.00154843, 0, 0.0346995, 0.0293831,
+ 0.0239779, 0.0184849, 0.012905, 0.0133686, 0.00943205, 0.00530731,
+ 0.00108283, 0, 0.00937699, 0.00689617, 0.00437921, 0.00182603,
+ 0, 0.00216168, 0.000431909, 0, 0, 0,
+ 0.0182273, 0.0184874, 0.018742, 0.0189907, 0.0137603, 0.0140486,
+ 0.0143348, 0.014619, 0.0149012, 0.012462, 0.0127637, 0.0131749,
+ 0.0137195, 0.0142671, 0.00858316, 0.00888649, 0.00919061, 0.00949552,
+ 0.00980122, 0.00658873, 0.00668349, 0.00677755, 0.00687091, 0.00696356,
+ 0, 0, 0, 0, 0.0026533, 0.00305218,
+ 0.00345251, 0.00385433, 0.00425764, 0.00128215, 0.00147873, 0.0016757,
+ 0.00187306, 0.00207081, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0.00312929, 0.00354451, 0.00396081, 0.00437819, 0, 0,
+ 0, 0, 0, 0.00283054, 0.00324669, 0.00366393,
+ 0.00408225, 0.00450167, 0.00320158, 0.00351594, 0.00383091, 0.00414651,
+ 0.00446272, 0.00477956, 0.0034087, 0.00361956, 0.0038307, 0.00404212,
+ 0.00425382, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0.00147984,
+ 0.00168904, 0.00189851, 0.00210825, 0)"
+          vdata_typ="(-1.8, -1.74, -1.68, -1.62, -1.56, -1.5,
+ -1.44, -1.38, -1.32, -1.26, -1.2, -1.14,
+ -1.08, -1.02, -0.96, -0.9, -0.84, -0.78,
+ -0.72, -0.66, -0.6, -0.54, -0.48, -0.42,
+ -0.36, -0.3, -0.24, -0.18, -0.12, -0.06,
+ 0, 0.06, 0.12, 0.18, 0.24, 0.3,
+ 0.36, 0.42, 0.48, 0.54, 0.6, 0.66,
+ 0.72, 0.78, 0.84, 0.9, 0.96, 1.02,
+ 1.08, 1.14, 1.2, 1.26, 1.32, 1.38,
+ 1.44, 1.5, 1.56, 1.62, 1.68, 1.74,
+ 1.8, 1.86, 1.92, 1.98, 2.04, 2.1,
+ 2.16, 2.22, 2.28, 2.34, 2.4, 2.46,
+ 2.52, 2.58, 2.64, 2.7, 2.76, 2.82,
+ 2.88, 2.94, 3, 3.06, 3.12, 3.18,
+ 3.24, 3.3, 3.36, 3.42, 3.48, 3.54,
+ 3.6)"
+          idata_typ="(-6.345, -5.918, -5.492, -5.066, -4.64, -4.214,
+ -3.788, -3.363, -2.937, -2.511, -2.086, -1.663,
+ -1.243, -0.8341, -0.4448, -0.196, -0.1389, -0.1177,
+ -0.1018, -0.08764, -0.075, -0.06428, -0.05584, -0.04952,
+ -0.04448, -0.0399, -0.03541, -0.03094, -0.02644, -0.02194,
+ -0.01743, -0.01301, -0.008738, -0.004612, -0.0006315, 0.003204,
+ 0.006895, 0.01044, 0.01383, 0.01707, 0.02014, 0.02303,
+ 0.02573, 0.02821, 0.03045, 0.03244, 0.0342, 0.03576,
+ 0.03718, 0.03853, 0.03986, 0.0412, 0.04257, 0.04398,
+ 0.04543, 0.04695, 0.04854, 0.0502, 0.05195, 0.05377,
+ 0.05569, 0.0577, 0.05975, 0.06183, 0.06393, 0.06606,
+ 0.06826, 0.07067, 0.07359, 0.0773, 0.08184, 0.08709,
+ 0.09294, 0.09942, 0.1074, 0.1257, 0.2032, 0.3338,
+ 0.4821, 0.6392, 0.7982, 0.9575, 1.116, 1.276,
+ 1.435, 1.595, 1.754, 1.914, 2.073, 2.233,
+ 2.392)"
+          tdata_0to1_min="(1.63161e-011, 2.2246e-011, 2.81759e-011, 3.41058e-011, 4.00356e-011, 4.59655e-011,
+ 5.18954e-011, 5.78253e-011, 6.37551e-011, 6.9685e-011, 7.56149e-011, 8.15448e-011,
+ 8.74746e-011, 9.34045e-011, 9.93344e-011, 1.05264e-010, 1.11194e-010, 1.17124e-010,
+ 1.23054e-010, 1.28984e-010, 1.34914e-010, 1.40843e-010, 1.46773e-010, 1.52703e-010,
+ 1.58633e-010, 1.64563e-010, 1.70493e-010, 1.76423e-010, 1.82353e-010, 1.88282e-010,
+ 1.94212e-010, 2.00142e-010, 2.06072e-010, 2.12002e-010, 2.17932e-010, 2.23862e-010,
+ 2.29792e-010, 2.35721e-010, 2.41651e-010, 2.47581e-010, 2.53511e-010, 2.59441e-010,
+ 2.65371e-010, 2.71301e-010, 2.77231e-010, 2.8316e-010, 2.8909e-010, 2.9502e-010,
+ 3.0095e-010, 3.0688e-010, 3.1281e-010, 3.1874e-010, 3.2467e-010, 3.30599e-010,
+ 3.36529e-010, 3.42459e-010, 3.48389e-010, 3.54319e-010, 3.60249e-010, 3.66179e-010,
+ 3.72109e-010, 3.78038e-010, 3.83968e-010, 3.89898e-010, 3.95828e-010, 4.01758e-010,
+ 4.07688e-010, 4.13618e-010, 4.19548e-010, 4.25477e-010, 4.31407e-010, 4.37337e-010,
+ 4.43267e-010, 4.49197e-010, 4.55127e-010, 4.61057e-010, 4.66987e-010, 4.72916e-010,
+ 4.78846e-010, 4.84776e-010, 4.90706e-010, 4.96636e-010, 5.02566e-010, 5.08496e-010,
+ 5.14426e-010, 5.20355e-010, 5.26285e-010, 5.32215e-010, 5.38145e-010, 5.44075e-010,
+ 5.50005e-010, 5.55935e-010, 5.61865e-010, 5.67794e-010, 5.73724e-010, 5.79654e-010,
+ 5.85584e-010, 5.91514e-010, 5.97444e-010, 6.03374e-010, 6.09304e-010, 6.15233e-010,
+ 6.21163e-010, 6.27093e-010, 6.33023e-010, 6.38953e-010, 6.44883e-010, 6.50813e-010,
+ 6.56743e-010, 6.62672e-010, 6.68602e-010, 6.74532e-010, 6.80462e-010, 6.86392e-010,
+ 6.92322e-010, 6.98252e-010, 7.04182e-010, 7.10111e-010, 7.16041e-010, 7.21971e-010,
+ 7.27901e-010, 7.33831e-010, 7.39761e-010, 7.45691e-010, 7.51621e-010, 7.5755e-010,
+ 7.6348e-010, 7.6941e-010, 7.7534e-010, 7.8127e-010, 7.872e-010, 7.9313e-010,
+ 7.9906e-010, 8.04989e-010, 8.10919e-010, 8.16849e-010, 8.22779e-010, 8.28709e-010,
+ 8.34639e-010, 8.40569e-010, 8.46499e-010, 8.52428e-010, 8.58358e-010, 8.64288e-010,
+ 8.70218e-010, 8.76148e-010, 8.82078e-010, 8.88008e-010, 8.93938e-010, 8.99867e-010,
+ 9.05797e-010, 9.11727e-010, 9.17657e-010, 9.23587e-010, 9.29517e-010, 9.35447e-010,
+ 9.41377e-010, 9.47306e-010, 9.53236e-010, 9.59166e-010, 9.65096e-010, 9.71026e-010,
+ 9.76956e-010, 9.82886e-010, 9.88816e-010, 9.94745e-010, 1.00068e-009, 1.00661e-009,
+ 1.01254e-009, 1.01846e-009, 1.02439e-009, 1.03032e-009, 1.03625e-009, 1.04218e-009,
+ 1.04811e-009, 1.05404e-009, 1.05997e-009, 1.0659e-009, 1.07183e-009, 1.07776e-009,
+ 1.08369e-009, 1.08962e-009, 1.09555e-009, 1.10148e-009, 1.10741e-009, 1.11334e-009,
+ 1.11927e-009, 1.1252e-009, 1.13113e-009, 1.13706e-009, 1.14299e-009, 1.14892e-009,
+ 1.15485e-009, 1.16078e-009, 1.16671e-009, 1.17264e-009, 1.17857e-009, 1.1845e-009,
+ 1.19043e-009, 1.19636e-009, 1.20229e-009, 1.20822e-009)"
+          kdata_0to1_min="(0, 0.00693597, 0.00734267, 0.00775038, 0.00815913, 0.00858505,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0.0149774, 0.0168403, 0.0186985, 0.0205519,
+ 0.0224006, 0.0240851, 0.0257124, 0.0534193, 0.0575498, 0.0616171,
+ 0.0656214, 0.069563, 0.102944, 0.109289, 0.1155, 0.121575,
+ 0.127512, 0.185885, 0.194014, 0.201885, 0.209487, 0.216904,
+ 0.262763, 0.270595, 0.278029, 0.284935, 0.291331, 0.389536,
+ 0.397239, 0.403807, 0.409531, 0.41272, 0.458302, 0.460574,
+ 0.460332, 0.45866, 0.456168, 0.521521, 0.519402, 0.516554,
+ 0.512182, 0.507981, 0.562714, 0.560143, 0.557616, 0.556013,
+ 0.55331, 0.659015, 0.662791, 0.666581, 0.669294, 0.672524,
+ 0.716442, 0.724711, 0.731962, 0.740509, 0.749691, 0.739752,
+ 0.749267, 0.759439, 0.770012, 0.780565, 0.791097, 0.79587,
+ 0.809271, 0.822809, 0.836161, 0.849325, 0.834494, 0.847778,
+ 0.862015, 0.876457, 0.891109, 0.864523, 0.877546, 0.890758,
+ 0.904235, 0.918949, 0.917735, 0.932302, 0.946993, 0.961955,
+ 0.977195, 0.924242, 0.935102, 0.946108, 0.957264, 0.968572,
+ 0.909004, 0.915836, 0.922722, 0.929662, 0.936656, 0.952113,
+ 0.960445, 0.968871, 0.977393, 0.986011, 0.960073, 0.966314,
+ 0.972606, 0.97895, 0.985348, 0.970999, 0.976042, 0.98112,
+ 0.986232, 0.991379, 0.972387, 0.975803, 0.979234, 0.98268,
+ 0.986141, 0.967094, 0.968918, 0.970746, 0.972578, 0.974414,
+ 0.973267, 0.97489, 0.976515, 0.978144, 0.979776, 0.98008,
+ 0.981606, 0.983135, 0.984771, 0.986428, 0.984285, 0.985785,
+ 0.987287, 0.988793, 0.990302, 0.982654, 0.983469, 0.984284,
+ 0.9851, 0.985918, 0.989565, 0.990614, 0.991664, 0.992715,
+ 0.993768, 0.993327, 0.994265, 0.995205, 0.996146, 0.997089,
+ 0.998032, 1, 1, 1, 1, 1,
+ 0.99667, 0.997028, 0.997387, 0.997745, 0.998104, 0.993811,
+ 0.993821, 0.99383, 0.99384, 0.993849, 0.998489, 0.998848,
+ 0.999207, 0.999566, 0.999926, 0.998882, 0.999149, 0.999417,
+ 0.999684, 0.999951, 1, 1)"
+          tdata_1to0_min="(7.19709e-011, 7.82209e-011, 8.44709e-011, 9.07209e-011, 9.69709e-011, 1.03221e-010,
+ 1.09471e-010, 1.15721e-010, 1.21971e-010, 1.28221e-010, 1.34471e-010, 1.40721e-010,
+ 1.46971e-010, 1.53221e-010, 1.59471e-010, 1.65721e-010, 1.71971e-010, 1.78221e-010,
+ 1.84471e-010, 1.90721e-010, 1.96971e-010, 2.03221e-010, 2.09471e-010, 2.15721e-010,
+ 2.21971e-010, 2.28221e-010, 2.34471e-010, 2.40721e-010, 2.46971e-010, 2.53221e-010,
+ 2.59471e-010, 2.65721e-010, 2.71971e-010, 2.78221e-010, 2.84471e-010, 2.90721e-010,
+ 2.96971e-010, 3.03221e-010, 3.09471e-010, 3.15721e-010, 3.21971e-010, 3.28221e-010,
+ 3.34471e-010, 3.40721e-010, 3.46971e-010, 3.53221e-010, 3.59471e-010, 3.65721e-010,
+ 3.71971e-010, 3.78221e-010, 3.84471e-010, 3.90721e-010, 3.96971e-010, 4.03221e-010,
+ 4.09471e-010, 4.15721e-010, 4.21971e-010, 4.28221e-010, 4.34471e-010, 4.40721e-010,
+ 4.46971e-010, 4.53221e-010, 4.59471e-010, 4.65721e-010, 4.71971e-010, 4.78221e-010,
+ 4.84471e-010, 4.90721e-010, 4.96971e-010, 5.03221e-010, 5.09471e-010, 5.15721e-010,
+ 5.21971e-010, 5.28221e-010, 5.34471e-010, 5.40721e-010, 5.46971e-010, 5.53221e-010,
+ 5.59471e-010, 5.65721e-010, 5.71971e-010, 5.78221e-010, 5.84471e-010, 5.90721e-010,
+ 5.96971e-010, 6.03221e-010, 6.09471e-010, 6.15721e-010, 6.21971e-010, 6.28221e-010,
+ 6.34471e-010, 6.40721e-010, 6.46971e-010, 6.53221e-010, 6.59471e-010, 6.65721e-010,
+ 6.71971e-010, 6.78221e-010, 6.84471e-010, 6.90721e-010, 6.96971e-010, 7.03221e-010,
+ 7.09471e-010, 7.15721e-010, 7.21971e-010, 7.28221e-010, 7.34471e-010, 7.40721e-010,
+ 7.46971e-010, 7.53221e-010, 7.59471e-010, 7.65721e-010, 7.71971e-010, 7.78221e-010,
+ 7.84471e-010, 7.90721e-010, 7.96971e-010, 8.03221e-010, 8.09471e-010, 8.15721e-010,
+ 8.21971e-010, 8.28221e-010, 8.34471e-010, 8.40721e-010, 8.46971e-010, 8.53221e-010,
+ 8.59471e-010, 8.65721e-010, 8.71971e-010, 8.78221e-010, 8.84471e-010, 8.90721e-010,
+ 8.96971e-010, 9.03221e-010, 9.09471e-010, 9.15721e-010, 9.21971e-010, 9.28221e-010,
+ 9.34471e-010, 9.40721e-010, 9.46971e-010, 9.53221e-010, 9.59471e-010, 9.65721e-010,
+ 9.71971e-010, 9.78221e-010, 9.84471e-010, 9.90721e-010, 9.96971e-010, 1.00322e-009,
+ 1.00947e-009, 1.01572e-009, 1.02197e-009, 1.02822e-009, 1.03447e-009, 1.04072e-009,
+ 1.04697e-009, 1.05322e-009, 1.05947e-009, 1.06572e-009, 1.07197e-009, 1.07822e-009,
+ 1.08447e-009, 1.09072e-009, 1.09697e-009, 1.10322e-009, 1.10947e-009, 1.11572e-009,
+ 1.12197e-009, 1.12822e-009, 1.13447e-009, 1.14072e-009, 1.14697e-009, 1.15322e-009,
+ 1.15947e-009, 1.16572e-009, 1.17197e-009, 1.17822e-009, 1.18447e-009, 1.19072e-009,
+ 1.19697e-009, 1.20322e-009, 1.20947e-009, 1.21572e-009, 1.22197e-009, 1.22822e-009,
+ 1.23447e-009, 1.24072e-009, 1.24697e-009, 1.25322e-009, 1.25947e-009, 1.26572e-009,
+ 1.27197e-009, 1.27822e-009, 1.28447e-009, 1.29072e-009, 1.29697e-009, 1.30322e-009,
+ 1.30947e-009, 1.31572e-009, 1.32197e-009, 1.32822e-009)"
+          kdata_1to0_min="(1, 0.969945, 0.967761, 0.965584, 0.963414, 0.961251,
+ 0.922663, 0.917876, 0.913122, 0.908402, 0.903714, 0.851047,
+ 0.843315, 0.835827, 0.828581, 0.821414, 0.777789, 0.768792,
+ 0.759918, 0.751166, 0.742532, 0.734016, 0.55307, 0.537138,
+ 0.52166, 0.506619, 0.491996, 0.366398, 0.350055, 0.334232,
+ 0.318906, 0.304052, 0.267484, 0.253148, 0.23932, 0.225815,
+ 0.212624, 0.239538, 0.228337, 0.217242, 0.206183, 0.204381,
+ 0.194033, 0.183877, 0.173777, 0.163736, 0.198952, 0.190664,
+ 0.182312, 0.1739, 0.165717, 0.170127, 0.16219, 0.154145,
+ 0.146131, 0.138011, 0.141711, 0.13341, 0.124857, 0.116071,
+ 0.107027, 0.153405, 0.145329, 0.136956, 0.128286, 0.11476,
+ 0.103503, 0.0919088, 0.0799865, 0.0670827, 0.0281211, 0.0117597,
+ 0, 0, 0, 0.0834382, 0.0701074, 0.0565091,
+ 0.0408893, 0.0245442, 0.0671925, 0.0543346, 0.0413051, 0.0277456,
+ 0.0127862, 0.00102775, 0, 0, 0, 0,
+ 0.0193647, 0.0104846, 0.00154843, 0, 0.0346995, 0.0293831,
+ 0.0239779, 0.0184849, 0.012905, 0.0133686, 0.00943205, 0.00530731,
+ 0.00108283, 0, 0.00937699, 0.00689617, 0.00437921, 0.00182603,
+ 0, 0.00216168, 0.000431909, 0, 0, 0,
+ 0.0182273, 0.0184874, 0.018742, 0.0189907, 0.0137603, 0.0140486,
+ 0.0143348, 0.014619, 0.0149012, 0.012462, 0.0127637, 0.0131749,
+ 0.0137195, 0.0142671, 0.00858316, 0.00888649, 0.00919061, 0.00949552,
+ 0.00980122, 0.00658873, 0.00668349, 0.00677755, 0.00687091, 0.00696356,
+ 0, 0, 0, 0, 0.0026533, 0.00305218,
+ 0.00345251, 0.00385433, 0.00425764, 0.00128215, 0.00147873, 0.0016757,
+ 0.00187306, 0.00207081, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0.00312929, 0.00354451, 0.00396081, 0.00437819, 0, 0,
+ 0, 0, 0, 0.00283054, 0.00324669, 0.00366393,
+ 0.00408225, 0.00450167, 0.00320158, 0.00351594, 0.00383091, 0.00414651,
+ 0.00446272, 0.00477956, 0.0034087, 0.00361956, 0.0038307, 0.00404212,
+ 0.00425382, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0.00147984,
+ 0.00168904, 0.00189851, 0.00210825, 0)"
+          vdata_min="(-1.8, -1.74, -1.68, -1.62, -1.56, -1.5,
+ -1.44, -1.38, -1.32, -1.26, -1.2, -1.14,
+ -1.08, -1.02, -0.96, -0.9, -0.84, -0.78,
+ -0.72, -0.66, -0.6, -0.54, -0.48, -0.42,
+ -0.36, -0.3, -0.24, -0.18, -0.12, -0.06,
+ 0, 0.06, 0.12, 0.18, 0.24, 0.3,
+ 0.36, 0.42, 0.48, 0.54, 0.6, 0.66,
+ 0.72, 0.78, 0.84, 0.9, 0.96, 1.02,
+ 1.08, 1.14, 1.2, 1.26, 1.32, 1.38,
+ 1.44, 1.5, 1.56, 1.62, 1.68, 1.74,
+ 1.8, 1.86, 1.92, 1.98, 2.04, 2.1,
+ 2.16, 2.22, 2.28, 2.34, 2.4, 2.46,
+ 2.52, 2.58, 2.64, 2.7, 2.76, 2.82,
+ 2.88, 2.94, 3, 3.06, 3.12, 3.18,
+ 3.24, 3.3, 3.36, 3.42, 3.48, 3.54,
+ 3.6)"
+          idata_min="(-6.345, -5.918, -5.492, -5.066, -4.64, -4.214,
+ -3.788, -3.363, -2.937, -2.511, -2.086, -1.663,
+ -1.243, -0.8341, -0.4448, -0.196, -0.1389, -0.1177,
+ -0.1018, -0.08764, -0.075, -0.06428, -0.05584, -0.04952,
+ -0.04448, -0.0399, -0.03541, -0.03094, -0.02644, -0.02194,
+ -0.01743, -0.01301, -0.008738, -0.004612, -0.0006315, 0.003204,
+ 0.006895, 0.01044, 0.01383, 0.01707, 0.02014, 0.02303,
+ 0.02573, 0.02821, 0.03045, 0.03244, 0.0342, 0.03576,
+ 0.03718, 0.03853, 0.03986, 0.0412, 0.04257, 0.04398,
+ 0.04543, 0.04695, 0.04854, 0.0502, 0.05195, 0.05377,
+ 0.05569, 0.0577, 0.05975, 0.06183, 0.06393, 0.06606,
+ 0.06826, 0.07067, 0.07359, 0.0773, 0.08184, 0.08709,
+ 0.09294, 0.09942, 0.1074, 0.1257, 0.2032, 0.3338,
+ 0.4821, 0.6392, 0.7982, 0.9575, 1.116, 1.276,
+ 1.435, 1.595, 1.754, 1.914, 2.073, 2.233,
+ 2.392)"
+          tdata_0to1_max="(1.63161e-011, 2.2246e-011, 2.81759e-011, 3.41058e-011, 4.00356e-011, 4.59655e-011,
+ 5.18954e-011, 5.78253e-011, 6.37551e-011, 6.9685e-011, 7.56149e-011, 8.15448e-011,
+ 8.74746e-011, 9.34045e-011, 9.93344e-011, 1.05264e-010, 1.11194e-010, 1.17124e-010,
+ 1.23054e-010, 1.28984e-010, 1.34914e-010, 1.40843e-010, 1.46773e-010, 1.52703e-010,
+ 1.58633e-010, 1.64563e-010, 1.70493e-010, 1.76423e-010, 1.82353e-010, 1.88282e-010,
+ 1.94212e-010, 2.00142e-010, 2.06072e-010, 2.12002e-010, 2.17932e-010, 2.23862e-010,
+ 2.29792e-010, 2.35721e-010, 2.41651e-010, 2.47581e-010, 2.53511e-010, 2.59441e-010,
+ 2.65371e-010, 2.71301e-010, 2.77231e-010, 2.8316e-010, 2.8909e-010, 2.9502e-010,
+ 3.0095e-010, 3.0688e-010, 3.1281e-010, 3.1874e-010, 3.2467e-010, 3.30599e-010,
+ 3.36529e-010, 3.42459e-010, 3.48389e-010, 3.54319e-010, 3.60249e-010, 3.66179e-010,
+ 3.72109e-010, 3.78038e-010, 3.83968e-010, 3.89898e-010, 3.95828e-010, 4.01758e-010,
+ 4.07688e-010, 4.13618e-010, 4.19548e-010, 4.25477e-010, 4.31407e-010, 4.37337e-010,
+ 4.43267e-010, 4.49197e-010, 4.55127e-010, 4.61057e-010, 4.66987e-010, 4.72916e-010,
+ 4.78846e-010, 4.84776e-010, 4.90706e-010, 4.96636e-010, 5.02566e-010, 5.08496e-010,
+ 5.14426e-010, 5.20355e-010, 5.26285e-010, 5.32215e-010, 5.38145e-010, 5.44075e-010,
+ 5.50005e-010, 5.55935e-010, 5.61865e-010, 5.67794e-010, 5.73724e-010, 5.79654e-010,
+ 5.85584e-010, 5.91514e-010, 5.97444e-010, 6.03374e-010, 6.09304e-010, 6.15233e-010,
+ 6.21163e-010, 6.27093e-010, 6.33023e-010, 6.38953e-010, 6.44883e-010, 6.50813e-010,
+ 6.56743e-010, 6.62672e-010, 6.68602e-010, 6.74532e-010, 6.80462e-010, 6.86392e-010,
+ 6.92322e-010, 6.98252e-010, 7.04182e-010, 7.10111e-010, 7.16041e-010, 7.21971e-010,
+ 7.27901e-010, 7.33831e-010, 7.39761e-010, 7.45691e-010, 7.51621e-010, 7.5755e-010,
+ 7.6348e-010, 7.6941e-010, 7.7534e-010, 7.8127e-010, 7.872e-010, 7.9313e-010,
+ 7.9906e-010, 8.04989e-010, 8.10919e-010, 8.16849e-010, 8.22779e-010, 8.28709e-010,
+ 8.34639e-010, 8.40569e-010, 8.46499e-010, 8.52428e-010, 8.58358e-010, 8.64288e-010,
+ 8.70218e-010, 8.76148e-010, 8.82078e-010, 8.88008e-010, 8.93938e-010, 8.99867e-010,
+ 9.05797e-010, 9.11727e-010, 9.17657e-010, 9.23587e-010, 9.29517e-010, 9.35447e-010,
+ 9.41377e-010, 9.47306e-010, 9.53236e-010, 9.59166e-010, 9.65096e-010, 9.71026e-010,
+ 9.76956e-010, 9.82886e-010, 9.88816e-010, 9.94745e-010, 1.00068e-009, 1.00661e-009,
+ 1.01254e-009, 1.01846e-009, 1.02439e-009, 1.03032e-009, 1.03625e-009, 1.04218e-009,
+ 1.04811e-009, 1.05404e-009, 1.05997e-009, 1.0659e-009, 1.07183e-009, 1.07776e-009,
+ 1.08369e-009, 1.08962e-009, 1.09555e-009, 1.10148e-009, 1.10741e-009, 1.11334e-009,
+ 1.11927e-009, 1.1252e-009, 1.13113e-009, 1.13706e-009, 1.14299e-009, 1.14892e-009,
+ 1.15485e-009, 1.16078e-009, 1.16671e-009, 1.17264e-009, 1.17857e-009, 1.1845e-009,
+ 1.19043e-009, 1.19636e-009, 1.20229e-009, 1.20822e-009)"
+          kdata_0to1_max="(0, 0.00693597, 0.00734267, 0.00775038, 0.00815913, 0.00858505,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0, 0, 0.0149774, 0.0168403, 0.0186985, 0.0205519,
+ 0.0224006, 0.0240851, 0.0257124, 0.0534193, 0.0575498, 0.0616171,
+ 0.0656214, 0.069563, 0.102944, 0.109289, 0.1155, 0.121575,
+ 0.127512, 0.185885, 0.194014, 0.201885, 0.209487, 0.216904,
+ 0.262763, 0.270595, 0.278029, 0.284935, 0.291331, 0.389536,
+ 0.397239, 0.403807, 0.409531, 0.41272, 0.458302, 0.460574,
+ 0.460332, 0.45866, 0.456168, 0.521521, 0.519402, 0.516554,
+ 0.512182, 0.507981, 0.562714, 0.560143, 0.557616, 0.556013,
+ 0.55331, 0.659015, 0.662791, 0.666581, 0.669294, 0.672524,
+ 0.716442, 0.724711, 0.731962, 0.740509, 0.749691, 0.739752,
+ 0.749267, 0.759439, 0.770012, 0.780565, 0.791097, 0.79587,
+ 0.809271, 0.822809, 0.836161, 0.849325, 0.834494, 0.847778,
+ 0.862015, 0.876457, 0.891109, 0.864523, 0.877546, 0.890758,
+ 0.904235, 0.918949, 0.917735, 0.932302, 0.946993, 0.961955,
+ 0.977195, 0.924242, 0.935102, 0.946108, 0.957264, 0.968572,
+ 0.909004, 0.915836, 0.922722, 0.929662, 0.936656, 0.952113,
+ 0.960445, 0.968871, 0.977393, 0.986011, 0.960073, 0.966314,
+ 0.972606, 0.97895, 0.985348, 0.970999, 0.976042, 0.98112,
+ 0.986232, 0.991379, 0.972387, 0.975803, 0.979234, 0.98268,
+ 0.986141, 0.967094, 0.968918, 0.970746, 0.972578, 0.974414,
+ 0.973267, 0.97489, 0.976515, 0.978144, 0.979776, 0.98008,
+ 0.981606, 0.983135, 0.984771, 0.986428, 0.984285, 0.985785,
+ 0.987287, 0.988793, 0.990302, 0.982654, 0.983469, 0.984284,
+ 0.9851, 0.985918, 0.989565, 0.990614, 0.991664, 0.992715,
+ 0.993768, 0.993327, 0.994265, 0.995205, 0.996146, 0.997089,
+ 0.998032, 1, 1, 1, 1, 1,
+ 0.99667, 0.997028, 0.997387, 0.997745, 0.998104, 0.993811,
+ 0.993821, 0.99383, 0.99384, 0.993849, 0.998489, 0.998848,
+ 0.999207, 0.999566, 0.999926, 0.998882, 0.999149, 0.999417,
+ 0.999684, 0.999951, 1, 1)"
+          tdata_1to0_max="(7.19709e-011, 7.82209e-011, 8.44709e-011, 9.07209e-011, 9.69709e-011, 1.03221e-010,
+ 1.09471e-010, 1.15721e-010, 1.21971e-010, 1.28221e-010, 1.34471e-010, 1.40721e-010,
+ 1.46971e-010, 1.53221e-010, 1.59471e-010, 1.65721e-010, 1.71971e-010, 1.78221e-010,
+ 1.84471e-010, 1.90721e-010, 1.96971e-010, 2.03221e-010, 2.09471e-010, 2.15721e-010,
+ 2.21971e-010, 2.28221e-010, 2.34471e-010, 2.40721e-010, 2.46971e-010, 2.53221e-010,
+ 2.59471e-010, 2.65721e-010, 2.71971e-010, 2.78221e-010, 2.84471e-010, 2.90721e-010,
+ 2.96971e-010, 3.03221e-010, 3.09471e-010, 3.15721e-010, 3.21971e-010, 3.28221e-010,
+ 3.34471e-010, 3.40721e-010, 3.46971e-010, 3.53221e-010, 3.59471e-010, 3.65721e-010,
+ 3.71971e-010, 3.78221e-010, 3.84471e-010, 3.90721e-010, 3.96971e-010, 4.03221e-010,
+ 4.09471e-010, 4.15721e-010, 4.21971e-010, 4.28221e-010, 4.34471e-010, 4.40721e-010,
+ 4.46971e-010, 4.53221e-010, 4.59471e-010, 4.65721e-010, 4.71971e-010, 4.78221e-010,
+ 4.84471e-010, 4.90721e-010, 4.96971e-010, 5.03221e-010, 5.09471e-010, 5.15721e-010,
+ 5.21971e-010, 5.28221e-010, 5.34471e-010, 5.40721e-010, 5.46971e-010, 5.53221e-010,
+ 5.59471e-010, 5.65721e-010, 5.71971e-010, 5.78221e-010, 5.84471e-010, 5.90721e-010,
+ 5.96971e-010, 6.03221e-010, 6.09471e-010, 6.15721e-010, 6.21971e-010, 6.28221e-010,
+ 6.34471e-010, 6.40721e-010, 6.46971e-010, 6.53221e-010, 6.59471e-010, 6.65721e-010,
+ 6.71971e-010, 6.78221e-010, 6.84471e-010, 6.90721e-010, 6.96971e-010, 7.03221e-010,
+ 7.09471e-010, 7.15721e-010, 7.21971e-010, 7.28221e-010, 7.34471e-010, 7.40721e-010,
+ 7.46971e-010, 7.53221e-010, 7.59471e-010, 7.65721e-010, 7.71971e-010, 7.78221e-010,
+ 7.84471e-010, 7.90721e-010, 7.96971e-010, 8.03221e-010, 8.09471e-010, 8.15721e-010,
+ 8.21971e-010, 8.28221e-010, 8.34471e-010, 8.40721e-010, 8.46971e-010, 8.53221e-010,
+ 8.59471e-010, 8.65721e-010, 8.71971e-010, 8.78221e-010, 8.84471e-010, 8.90721e-010,
+ 8.96971e-010, 9.03221e-010, 9.09471e-010, 9.15721e-010, 9.21971e-010, 9.28221e-010,
+ 9.34471e-010, 9.40721e-010, 9.46971e-010, 9.53221e-010, 9.59471e-010, 9.65721e-010,
+ 9.71971e-010, 9.78221e-010, 9.84471e-010, 9.90721e-010, 9.96971e-010, 1.00322e-009,
+ 1.00947e-009, 1.01572e-009, 1.02197e-009, 1.02822e-009, 1.03447e-009, 1.04072e-009,
+ 1.04697e-009, 1.05322e-009, 1.05947e-009, 1.06572e-009, 1.07197e-009, 1.07822e-009,
+ 1.08447e-009, 1.09072e-009, 1.09697e-009, 1.10322e-009, 1.10947e-009, 1.11572e-009,
+ 1.12197e-009, 1.12822e-009, 1.13447e-009, 1.14072e-009, 1.14697e-009, 1.15322e-009,
+ 1.15947e-009, 1.16572e-009, 1.17197e-009, 1.17822e-009, 1.18447e-009, 1.19072e-009,
+ 1.19697e-009, 1.20322e-009, 1.20947e-009, 1.21572e-009, 1.22197e-009, 1.22822e-009,
+ 1.23447e-009, 1.24072e-009, 1.24697e-009, 1.25322e-009, 1.25947e-009, 1.26572e-009,
+ 1.27197e-009, 1.27822e-009, 1.28447e-009, 1.29072e-009, 1.29697e-009, 1.30322e-009,
+ 1.30947e-009, 1.31572e-009, 1.32197e-009, 1.32822e-009)"
+          kdata_1to0_max="(1, 0.969945, 0.967761, 0.965584, 0.963414, 0.961251,
+ 0.922663, 0.917876, 0.913122, 0.908402, 0.903714, 0.851047,
+ 0.843315, 0.835827, 0.828581, 0.821414, 0.777789, 0.768792,
+ 0.759918, 0.751166, 0.742532, 0.734016, 0.55307, 0.537138,
+ 0.52166, 0.506619, 0.491996, 0.366398, 0.350055, 0.334232,
+ 0.318906, 0.304052, 0.267484, 0.253148, 0.23932, 0.225815,
+ 0.212624, 0.239538, 0.228337, 0.217242, 0.206183, 0.204381,
+ 0.194033, 0.183877, 0.173777, 0.163736, 0.198952, 0.190664,
+ 0.182312, 0.1739, 0.165717, 0.170127, 0.16219, 0.154145,
+ 0.146131, 0.138011, 0.141711, 0.13341, 0.124857, 0.116071,
+ 0.107027, 0.153405, 0.145329, 0.136956, 0.128286, 0.11476,
+ 0.103503, 0.0919088, 0.0799865, 0.0670827, 0.0281211, 0.0117597,
+ 0, 0, 0, 0.0834382, 0.0701074, 0.0565091,
+ 0.0408893, 0.0245442, 0.0671925, 0.0543346, 0.0413051, 0.0277456,
+ 0.0127862, 0.00102775, 0, 0, 0, 0,
+ 0.0193647, 0.0104846, 0.00154843, 0, 0.0346995, 0.0293831,
+ 0.0239779, 0.0184849, 0.012905, 0.0133686, 0.00943205, 0.00530731,
+ 0.00108283, 0, 0.00937699, 0.00689617, 0.00437921, 0.00182603,
+ 0, 0.00216168, 0.000431909, 0, 0, 0,
+ 0.0182273, 0.0184874, 0.018742, 0.0189907, 0.0137603, 0.0140486,
+ 0.0143348, 0.014619, 0.0149012, 0.012462, 0.0127637, 0.0131749,
+ 0.0137195, 0.0142671, 0.00858316, 0.00888649, 0.00919061, 0.00949552,
+ 0.00980122, 0.00658873, 0.00668349, 0.00677755, 0.00687091, 0.00696356,
+ 0, 0, 0, 0, 0.0026533, 0.00305218,
+ 0.00345251, 0.00385433, 0.00425764, 0.00128215, 0.00147873, 0.0016757,
+ 0.00187306, 0.00207081, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0,
+ 0.00312929, 0.00354451, 0.00396081, 0.00437819, 0, 0,
+ 0, 0, 0, 0.00283054, 0.00324669, 0.00366393,
+ 0.00408225, 0.00450167, 0.00320158, 0.00351594, 0.00383091, 0.00414651,
+ 0.00446272, 0.00477956, 0.0034087, 0.00361956, 0.0038307, 0.00404212,
+ 0.00425382, 0, 0, 0, 0, 0,
+ 0, 0, 0, 0, 0, 0.00147984,
+ 0.00168904, 0.00189851, 0.00210825, 0)"
+          vdata_max="(-1.8, -1.74, -1.68, -1.62, -1.56, -1.5,
+ -1.44, -1.38, -1.32, -1.26, -1.2, -1.14,
+ -1.08, -1.02, -0.96, -0.9, -0.84, -0.78,
+ -0.72, -0.66, -0.6, -0.54, -0.48, -0.42,
+ -0.36, -0.3, -0.24, -0.18, -0.12, -0.06,
+ 0, 0.06, 0.12, 0.18, 0.24, 0.3,
+ 0.36, 0.42, 0.48, 0.54, 0.6, 0.66,
+ 0.72, 0.78, 0.84, 0.9, 0.96, 1.02,
+ 1.08, 1.14, 1.2, 1.26, 1.32, 1.38,
+ 1.44, 1.5, 1.56, 1.62, 1.68, 1.74,
+ 1.8, 1.86, 1.92, 1.98, 2.04, 2.1,
+ 2.16, 2.22, 2.28, 2.34, 2.4, 2.46,
+ 2.52, 2.58, 2.64, 2.7, 2.76, 2.82,
+ 2.88, 2.94, 3, 3.06, 3.12, 3.18,
+ 3.24, 3.3, 3.36, 3.42, 3.48, 3.54,
+ 3.6)"
+          idata_max="(-6.345, -5.918, -5.492, -5.066, -4.64, -4.214,
+ -3.788, -3.363, -2.937, -2.511, -2.086, -1.663,
+ -1.243, -0.8341, -0.4448, -0.196, -0.1389, -0.1177,
+ -0.1018, -0.08764, -0.075, -0.06428, -0.05584, -0.04952,
+ -0.04448, -0.0399, -0.03541, -0.03094, -0.02644, -0.02194,
+ -0.01743, -0.01301, -0.008738, -0.004612, -0.0006315, 0.003204,
+ 0.006895, 0.01044, 0.01383, 0.01707, 0.02014, 0.02303,
+ 0.02573, 0.02821, 0.03045, 0.03244, 0.0342, 0.03576,
+ 0.03718, 0.03853, 0.03986, 0.0412, 0.04257, 0.04398,
+ 0.04543, 0.04695, 0.04854, 0.0502, 0.05195, 0.05377,
+ 0.05569, 0.0577, 0.05975, 0.06183, 0.06393, 0.06606,
+ 0.06826, 0.07067, 0.07359, 0.0773, 0.08184, 0.08709,
+ 0.09294, 0.09942, 0.1074, 0.1257, 0.2032, 0.3338,
+ 0.4821, 0.6392, 0.7982, 0.9575, 1.116, 1.276,
+ 1.435, 1.595, 1.754, 1.914, 2.073, 2.233,
+ 2.392)"
+ PORT: a_PdRef
+       a_signal
+       d_pulldown_control


*IBIS Pullup tables
Y_PullUp ibis_ktiv(icx_behavioral)
+ GENERIC: corner="ibis_typ"
+          tdata_0to1_typ="(7.19709e-011, 7.82209e-011, 8.44709e-011, 9.07209e-011, 9.69709e-011, 1.03221e-010,
+ 1.09471e-010, 1.15721e-010, 1.21971e-010, 1.28221e-010, 1.34471e-010, 1.40721e-010,
+ 1.46971e-010, 1.53221e-010, 1.59471e-010, 1.65721e-010, 1.71971e-010, 1.78221e-010,
+ 1.84471e-010, 1.90721e-010, 1.96971e-010, 2.03221e-010, 2.09471e-010, 2.15721e-010,
+ 2.21971e-010, 2.28221e-010, 2.34471e-010, 2.40721e-010, 2.46971e-010, 2.53221e-010,
+ 2.59471e-010, 2.65721e-010, 2.71971e-010, 2.78221e-010, 2.84471e-010, 2.90721e-010,
+ 2.96971e-010, 3.03221e-010, 3.09471e-010, 3.15721e-010, 3.21971e-010, 3.28221e-010,
+ 3.34471e-010, 3.40721e-010, 3.46971e-010, 3.53221e-010, 3.59471e-010, 3.65721e-010,
+ 3.71971e-010, 3.78221e-010, 3.84471e-010, 3.90721e-010, 3.96971e-010, 4.03221e-010,
+ 4.09471e-010, 4.15721e-010, 4.21971e-010, 4.28221e-010, 4.34471e-010, 4.40721e-010,
+ 4.46971e-010, 4.53221e-010, 4.59471e-010, 4.65721e-010, 4.71971e-010, 4.78221e-010,
+ 4.84471e-010, 4.90721e-010, 4.96971e-010, 5.03221e-010, 5.09471e-010, 5.15721e-010,
+ 5.21971e-010, 5.28221e-010, 5.34471e-010, 5.40721e-010, 5.46971e-010, 5.53221e-010,
+ 5.59471e-010, 5.65721e-010, 5.71971e-010, 5.78221e-010, 5.84471e-010, 5.90721e-010,
+ 5.96971e-010, 6.03221e-010, 6.09471e-010, 6.15721e-010, 6.21971e-010, 6.28221e-010,
+ 6.34471e-010, 6.40721e-010, 6.46971e-010, 6.53221e-010, 6.59471e-010, 6.65721e-010,
+ 6.71971e-010, 6.78221e-010, 6.84471e-010, 6.90721e-010, 6.96971e-010, 7.03221e-010,
+ 7.09471e-010, 7.15721e-010, 7.21971e-010, 7.28221e-010, 7.34471e-010, 7.40721e-010,
+ 7.46971e-010, 7.53221e-010, 7.59471e-010, 7.65721e-010, 7.71971e-010, 7.78221e-010,
+ 7.84471e-010, 7.90721e-010, 7.96971e-010, 8.03221e-010, 8.09471e-010, 8.15721e-010,
+ 8.21971e-010, 8.28221e-010, 8.34471e-010, 8.40721e-010, 8.46971e-010, 8.53221e-010,
+ 8.59471e-010, 8.65721e-010, 8.71971e-010, 8.78221e-010, 8.84471e-010, 8.90721e-010,
+ 8.96971e-010, 9.03221e-010, 9.09471e-010, 9.15721e-010, 9.21971e-010, 9.28221e-010,
+ 9.34471e-010, 9.40721e-010, 9.46971e-010, 9.53221e-010, 9.59471e-010, 9.65721e-010,
+ 9.71971e-010, 9.78221e-010, 9.84471e-010, 9.90721e-010, 9.96971e-010, 1.00322e-009,
+ 1.00947e-009, 1.01572e-009, 1.02197e-009, 1.02822e-009, 1.03447e-009, 1.04072e-009,
+ 1.04697e-009, 1.05322e-009, 1.05947e-009, 1.06572e-009, 1.07197e-009, 1.07822e-009,
+ 1.08447e-009, 1.09072e-009, 1.09697e-009, 1.10322e-009, 1.10947e-009, 1.11572e-009,
+ 1.12197e-009, 1.12822e-009, 1.13447e-009, 1.14072e-009, 1.14697e-009, 1.15322e-009,
+ 1.15947e-009, 1.16572e-009, 1.17197e-009, 1.17822e-009, 1.18447e-009, 1.19072e-009,
+ 1.19697e-009, 1.20322e-009, 1.20947e-009, 1.21572e-009, 1.22197e-009, 1.22822e-009,
+ 1.23447e-009, 1.24072e-009, 1.24697e-009, 1.25322e-009, 1.25947e-009, 1.26572e-009,
+ 1.27197e-009, 1.27822e-009, 1.28447e-009, 1.29072e-009, 1.29697e-009, 1.30322e-009,
+ 1.30947e-009, 1.31572e-009, 1.32197e-009, 1.32822e-009)"
+          kdata_0to1_typ="(0, 0.00144844, 0.00161591, 0.00178283, 0.00194921, 0.00211506,
+ 0.0087038, 0.00937234, 0.0100361, 0.0106951, 0.0113493, 0.0221732,
+ 0.0235462, 0.0248913, 0.0262091, 0.027512, 0.0384896, 0.040387,
+ 0.0422566, 0.0440992, 0.0459152, 0.0477052, 0.0909226, 0.0947716,
+ 0.0985008, 0.102115, 0.10562, 0.151672, 0.156561, 0.161263,
+ 0.165788, 0.170143, 0.231451, 0.237879, 0.244041, 0.249991,
+ 0.255738, 0.306646, 0.314487, 0.322133, 0.329544, 0.346723,
+ 0.354268, 0.361647, 0.368849, 0.375871, 0.436727, 0.446473,
+ 0.456075, 0.465528, 0.47489, 0.508024, 0.518296, 0.528421,
+ 0.538431, 0.548284, 0.578952, 0.589365, 0.599555, 0.609511,
+ 0.619187, 0.661993, 0.673295, 0.684356, 0.695153, 0.695174,
+ 0.703634, 0.711667, 0.719248, 0.725866, 0.705895, 0.708557,
+ 0.710598, 0.711564, 0.710588, 0.813801, 0.819259, 0.824199,
+ 0.827163, 0.82912, 0.854347, 0.858385, 0.861996, 0.865003,
+ 0.86646, 0.82184, 0.821897, 0.821674, 0.821592, 0.821429,
+ 0.86842, 0.871631, 0.874676, 0.877554, 0.928498, 0.936229,
+ 0.943903, 0.951517, 0.95907, 0.902802, 0.908617, 0.914903,
+ 0.921194, 0.927466, 0.912617, 0.919099, 0.925592, 0.932094,
+ 0.938605, 0.915914, 0.921739, 0.928803, 0.935927, 0.943095,
+ 0.982139, 0.992066, 1, 1, 0.970056, 0.977633,
+ 0.985279, 0.992996, 1, 0.981505, 0.988024, 0.995008,
+ 1, 1, 0.97652, 0.981778, 0.987072, 0.992403,
+ 0.997772, 0.989569, 0.994141, 0.99874, 1, 1,
+ 0.958503, 0.959695, 0.960888, 0.961952, 0.984313, 0.987439,
+ 0.99058, 0.993734, 0.996902, 0.986424, 0.988754, 0.991091,
+ 0.993435, 0.995786, 0.984205, 0.985709, 0.987216, 0.988726,
+ 0.990238, 0.991754, 0.993272, 0.994792, 0.996316, 0.997843,
+ 0.997771, 0.99948, 1, 1, 0.978729, 0.978557,
+ 0.978385, 0.978213, 0.978042, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 0.984196, 0.983159, 0.982125, 0.981093, 0.980062,
+ 0.991678, 0.991678, 0.991678, 0.991678, 0.991678, 1,
+ 1, 1, 1, 1)"
+          tdata_1to0_typ="(1.63161e-011, 2.2246e-011, 2.81759e-011, 3.41058e-011, 4.00356e-011, 4.59655e-011,
+ 5.18954e-011, 5.78253e-011, 6.37551e-011, 6.9685e-011, 7.56149e-011, 8.15448e-011,
+ 8.74746e-011, 9.34045e-011, 9.93344e-011, 1.05264e-010, 1.11194e-010, 1.17124e-010,
+ 1.23054e-010, 1.28984e-010, 1.34914e-010, 1.40843e-010, 1.46773e-010, 1.52703e-010,
+ 1.58633e-010, 1.64563e-010, 1.70493e-010, 1.76423e-010, 1.82353e-010, 1.88282e-010,
+ 1.94212e-010, 2.00142e-010, 2.06072e-010, 2.12002e-010, 2.17932e-010, 2.23862e-010,
+ 2.29792e-010, 2.35721e-010, 2.41651e-010, 2.47581e-010, 2.53511e-010, 2.59441e-010,
+ 2.65371e-010, 2.71301e-010, 2.77231e-010, 2.8316e-010, 2.8909e-010, 2.9502e-010,
+ 3.0095e-010, 3.0688e-010, 3.1281e-010, 3.1874e-010, 3.2467e-010, 3.30599e-010,
+ 3.36529e-010, 3.42459e-010, 3.48389e-010, 3.54319e-010, 3.60249e-010, 3.66179e-010,
+ 3.72109e-010, 3.78038e-010, 3.83968e-010, 3.89898e-010, 3.95828e-010, 4.01758e-010,
+ 4.07688e-010, 4.13618e-010, 4.19548e-010, 4.25477e-010, 4.31407e-010, 4.37337e-010,
+ 4.43267e-010, 4.49197e-010, 4.55127e-010, 4.61057e-010, 4.66987e-010, 4.72916e-010,
+ 4.78846e-010, 4.84776e-010, 4.90706e-010, 4.96636e-010, 5.02566e-010, 5.08496e-010,
+ 5.14426e-010, 5.20355e-010, 5.26285e-010, 5.32215e-010, 5.38145e-010, 5.44075e-010,
+ 5.50005e-010, 5.55935e-010, 5.61865e-010, 5.67794e-010, 5.73724e-010, 5.79654e-010,
+ 5.85584e-010, 5.91514e-010, 5.97444e-010, 6.03374e-010, 6.09304e-010, 6.15233e-010,
+ 6.21163e-010, 6.27093e-010, 6.33023e-010, 6.38953e-010, 6.44883e-010, 6.50813e-010,
+ 6.56743e-010, 6.62672e-010, 6.68602e-010, 6.74532e-010, 6.80462e-010, 6.86392e-010,
+ 6.92322e-010, 6.98252e-010, 7.04182e-010, 7.10111e-010, 7.16041e-010, 7.21971e-010,
+ 7.27901e-010, 7.33831e-010, 7.39761e-010, 7.45691e-010, 7.51621e-010, 7.5755e-010,
+ 7.6348e-010, 7.6941e-010, 7.7534e-010, 7.8127e-010, 7.872e-010, 7.9313e-010,
+ 7.9906e-010, 8.04989e-010, 8.10919e-010, 8.16849e-010, 8.22779e-010, 8.28709e-010,
+ 8.34639e-010, 8.40569e-010, 8.46499e-010, 8.52428e-010, 8.58358e-010, 8.64288e-010,
+ 8.70218e-010, 8.76148e-010, 8.82078e-010, 8.88008e-010, 8.93938e-010, 8.99867e-010,
+ 9.05797e-010, 9.11727e-010, 9.17657e-010, 9.23587e-010, 9.29517e-010, 9.35447e-010,
+ 9.41377e-010, 9.47306e-010, 9.53236e-010, 9.59166e-010, 9.65096e-010, 9.71026e-010,
+ 9.76956e-010, 9.82886e-010, 9.88816e-010, 9.94745e-010, 1.00068e-009, 1.00661e-009,
+ 1.01254e-009, 1.01846e-009, 1.02439e-009, 1.03032e-009, 1.03625e-009, 1.04218e-009,
+ 1.04811e-009, 1.05404e-009, 1.05997e-009, 1.0659e-009, 1.07183e-009, 1.07776e-009,
+ 1.08369e-009, 1.08962e-009, 1.09555e-009, 1.10148e-009, 1.10741e-009, 1.11334e-009,
+ 1.11927e-009, 1.1252e-009, 1.13113e-009, 1.13706e-009, 1.14299e-009, 1.14892e-009,
+ 1.15485e-009, 1.16078e-009, 1.16671e-009, 1.17264e-009, 1.17857e-009, 1.1845e-009,
+ 1.19043e-009, 1.19636e-009, 1.20229e-009, 1.20822e-009)"
+          kdata_1to0_typ="(1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 0.944958, 0.941817, 0.939014,
+ 0.936329, 0.933652, 0.928097, 0.926197, 0.924296, 0.922394,
+ 0.920489, 0.918327, 0.916081, 0.742328, 0.734287, 0.726279,
+ 0.718306, 0.710366, 0.5818, 0.572814, 0.563786, 0.554718,
+ 0.545614, 0.432759, 0.422287, 0.411632, 0.400804, 0.390031,
+ 0.357675, 0.345405, 0.33285, 0.319786, 0.306318, 0.299028,
+ 0.281999, 0.263834, 0.245179, 0.224, 0.21373, 0.19043,
+ 0.164822, 0.138767, 0.11283, 0.168453, 0.142421, 0.11653,
+ 0.0898447, 0.064093, 0.12499, 0.101151, 0.0779349, 0.0556811,
+ 0.0329568, 0.116942, 0.0977118, 0.0785584, 0.0587776, 0.0393621,
+ 0.100619, 0.0856291, 0.0698708, 0.0543328, 0.0388455, 0.0738995,
+ 0.0617298, 0.0492707, 0.0366203, 0.0238299, 0.0109021, 0.0561065,
+ 0.0467763, 0.0372812, 0.0274446, 0.0172799, 0.0457196, 0.0381295,
+ 0.0304268, 0.0225745, 0.0145697, 0.0383468, 0.0325389, 0.0266255,
+ 0.0206042, 0.0144643, 0.0365308, 0.0322321, 0.0277894, 0.0232542,
+ 0.0186239, 0.028672, 0.025203, 0.0216809, 0.0181047, 0.0144733,
+ 0.0148853, 0.0116153, 0.00831567, 0.00498609, 0.0016262, 0.0188761,
+ 0.0170186, 0.015139, 0.0132368, 0.0113117, 0.0155086, 0.0140556,
+ 0.0125899, 0.0111111, 0.00961925, 0.0139533, 0.0129102, 0.0118597,
+ 0.0108016, 0.00973602, 0.0114324, 0.0105801, 0.00972376, 0.00886338,
+ 0.00799891, 0.00901914, 0.00830074, 0.00758063, 0.0068588, 0.00613525,
+ 0.00561266, 0.00490209, 0.00419006, 0.00347656, 0.00276158, 0.00173159,
+ 0.000988725, 0.000244458, 0, 0, 0.00391781, 0.00364127,
+ 0.00336415, 0.00308644, 0.00280814, 0.00360153, 0.003408, 0.00321424,
+ 0.00302027, 0.00282607, 0.00282379, 0.00264561, 0.00246717, 0.00228846,
+ 0.00210949, 0.00204093, 0.00187022, 0.00169929, 0.00152814, 0.00135675,
+ 0.00118514, 0.00121595, 0.00106019, 0.000904174, 0.000747895, 0.000591352,
+ 0.00127719, 0.00118284, 0.00108844, 0.000993996, 0.000899505, 0.000727513,
+ 0.000625664, 0.000523821, 0.000421982, 0.000320148, 0.000293503, 0.000198808,
+ 0.000104067, 9.27975e-006, 0, 0.0004531, 0.000407536, 0.000361956,
+ 0.000316359, 0.000270744, 0.000225112, 0)"
+          vdata_typ="(-1.8, -1.74, -1.68, -1.62, -1.56, -1.5,
+ -1.44, -1.38, -1.32, -1.26, -1.2, -1.14,
+ -1.08, -1.02, -0.96, -0.9, -0.84, -0.78,
+ -0.72, -0.66, -0.6, -0.54, -0.48, -0.42,
+ -0.36, -0.3, -0.24, -0.18, -0.12, -0.06,
+ 0, 0.06, 0.12, 0.18, 0.24, 0.3,
+ 0.36, 0.42, 0.48, 0.54, 0.6, 0.66,
+ 0.72, 0.78, 0.84, 0.9, 0.96, 1.02,
+ 1.08, 1.14, 1.2, 1.26, 1.32, 1.38,
+ 1.44, 1.5, 1.56, 1.62, 1.68, 1.74,
+ 1.8, 1.86, 1.92, 1.98, 2.04, 2.1,
+ 2.16, 2.22, 2.28, 2.34, 2.4, 2.46,
+ 2.52, 2.58, 2.64, 2.7, 2.76, 2.82,
+ 2.88, 2.94, 3, 3.06, 3.12, 3.18,
+ 3.24, 3.3, 3.36, 3.42, 3.48, 3.54,
+ 3.6)"
+          idata_typ="(-2.394, -2.235, -2.075, -1.915, -1.756, -1.596,
+ -1.437, -1.277, -1.118, -0.9586, -0.7993, -0.6403,
+ -0.4841, -0.3375, -0.2096, -0.1333, -0.1135, -0.1032,
+ -0.09427, -0.08574, -0.07761, -0.06996, -0.06286, -0.05631,
+ -0.05017, -0.04422, -0.03837, -0.03258, -0.02687, -0.02127,
+ -0.01578, -0.01053, -0.005574, -0.0009032, 0.003482, 0.007583,
+ 0.0114, 0.01494, 0.0182, 0.02119, 0.0239, 0.02632,
+ 0.02844, 0.03027, 0.03189, 0.03338, 0.03481, 0.0362,
+ 0.03759, 0.03898, 0.04039, 0.04181, 0.04324, 0.0447,
+ 0.04617, 0.04766, 0.04918, 0.05073, 0.0523, 0.0539,
+ 0.05554, 0.05721, 0.05887, 0.06051, 0.06215, 0.06379,
+ 0.06553, 0.06774, 0.07132, 0.07727, 0.08581, 0.09653,
+ 0.109, 0.1233, 0.143, 0.1988, 0.4466, 0.8356,
+ 1.244, 1.664, 2.088, 2.513, 2.938, 3.364,
+ 3.79, 4.216, 4.641, 5.067, 5.493, 5.919,
+ 6.346)"
+          tdata_0to1_min="(7.19709e-011, 7.82209e-011, 8.44709e-011, 9.07209e-011, 9.69709e-011, 1.03221e-010,
+ 1.09471e-010, 1.15721e-010, 1.21971e-010, 1.28221e-010, 1.34471e-010, 1.40721e-010,
+ 1.46971e-010, 1.53221e-010, 1.59471e-010, 1.65721e-010, 1.71971e-010, 1.78221e-010,
+ 1.84471e-010, 1.90721e-010, 1.96971e-010, 2.03221e-010, 2.09471e-010, 2.15721e-010,
+ 2.21971e-010, 2.28221e-010, 2.34471e-010, 2.40721e-010, 2.46971e-010, 2.53221e-010,
+ 2.59471e-010, 2.65721e-010, 2.71971e-010, 2.78221e-010, 2.84471e-010, 2.90721e-010,
+ 2.96971e-010, 3.03221e-010, 3.09471e-010, 3.15721e-010, 3.21971e-010, 3.28221e-010,
+ 3.34471e-010, 3.40721e-010, 3.46971e-010, 3.53221e-010, 3.59471e-010, 3.65721e-010,
+ 3.71971e-010, 3.78221e-010, 3.84471e-010, 3.90721e-010, 3.96971e-010, 4.03221e-010,
+ 4.09471e-010, 4.15721e-010, 4.21971e-010, 4.28221e-010, 4.34471e-010, 4.40721e-010,
+ 4.46971e-010, 4.53221e-010, 4.59471e-010, 4.65721e-010, 4.71971e-010, 4.78221e-010,
+ 4.84471e-010, 4.90721e-010, 4.96971e-010, 5.03221e-010, 5.09471e-010, 5.15721e-010,
+ 5.21971e-010, 5.28221e-010, 5.34471e-010, 5.40721e-010, 5.46971e-010, 5.53221e-010,
+ 5.59471e-010, 5.65721e-010, 5.71971e-010, 5.78221e-010, 5.84471e-010, 5.90721e-010,
+ 5.96971e-010, 6.03221e-010, 6.09471e-010, 6.15721e-010, 6.21971e-010, 6.28221e-010,
+ 6.34471e-010, 6.40721e-010, 6.46971e-010, 6.53221e-010, 6.59471e-010, 6.65721e-010,
+ 6.71971e-010, 6.78221e-010, 6.84471e-010, 6.90721e-010, 6.96971e-010, 7.03221e-010,
+ 7.09471e-010, 7.15721e-010, 7.21971e-010, 7.28221e-010, 7.34471e-010, 7.40721e-010,
+ 7.46971e-010, 7.53221e-010, 7.59471e-010, 7.65721e-010, 7.71971e-010, 7.78221e-010,
+ 7.84471e-010, 7.90721e-010, 7.96971e-010, 8.03221e-010, 8.09471e-010, 8.15721e-010,
+ 8.21971e-010, 8.28221e-010, 8.34471e-010, 8.40721e-010, 8.46971e-010, 8.53221e-010,
+ 8.59471e-010, 8.65721e-010, 8.71971e-010, 8.78221e-010, 8.84471e-010, 8.90721e-010,
+ 8.96971e-010, 9.03221e-010, 9.09471e-010, 9.15721e-010, 9.21971e-010, 9.28221e-010,
+ 9.34471e-010, 9.40721e-010, 9.46971e-010, 9.53221e-010, 9.59471e-010, 9.65721e-010,
+ 9.71971e-010, 9.78221e-010, 9.84471e-010, 9.90721e-010, 9.96971e-010, 1.00322e-009,
+ 1.00947e-009, 1.01572e-009, 1.02197e-009, 1.02822e-009, 1.03447e-009, 1.04072e-009,
+ 1.04697e-009, 1.05322e-009, 1.05947e-009, 1.06572e-009, 1.07197e-009, 1.07822e-009,
+ 1.08447e-009, 1.09072e-009, 1.09697e-009, 1.10322e-009, 1.10947e-009, 1.11572e-009,
+ 1.12197e-009, 1.12822e-009, 1.13447e-009, 1.14072e-009, 1.14697e-009, 1.15322e-009,
+ 1.15947e-009, 1.16572e-009, 1.17197e-009, 1.17822e-009, 1.18447e-009, 1.19072e-009,
+ 1.19697e-009, 1.20322e-009, 1.20947e-009, 1.21572e-009, 1.22197e-009, 1.22822e-009,
+ 1.23447e-009, 1.24072e-009, 1.24697e-009, 1.25322e-009, 1.25947e-009, 1.26572e-009,
+ 1.27197e-009, 1.27822e-009, 1.28447e-009, 1.29072e-009, 1.29697e-009, 1.30322e-009,
+ 1.30947e-009, 1.31572e-009, 1.32197e-009, 1.32822e-009)"
+          kdata_0to1_min="(0, 0.00144844, 0.00161591, 0.00178283, 0.00194921, 0.00211506,
+ 0.0087038, 0.00937234, 0.0100361, 0.0106951, 0.0113493, 0.0221732,
+ 0.0235462, 0.0248913, 0.0262091, 0.027512, 0.0384896, 0.040387,
+ 0.0422566, 0.0440992, 0.0459152, 0.0477052, 0.0909226, 0.0947716,
+ 0.0985008, 0.102115, 0.10562, 0.151672, 0.156561, 0.161263,
+ 0.165788, 0.170143, 0.231451, 0.237879, 0.244041, 0.249991,
+ 0.255738, 0.306646, 0.314487, 0.322133, 0.329544, 0.346723,
+ 0.354268, 0.361647, 0.368849, 0.375871, 0.436727, 0.446473,
+ 0.456075, 0.465528, 0.47489, 0.508024, 0.518296, 0.528421,
+ 0.538431, 0.548284, 0.578952, 0.589365, 0.599555, 0.609511,
+ 0.619187, 0.661993, 0.673295, 0.684356, 0.695153, 0.695174,
+ 0.703634, 0.711667, 0.719248, 0.725866, 0.705895, 0.708557,
+ 0.710598, 0.711564, 0.710588, 0.813801, 0.819259, 0.824199,
+ 0.827163, 0.82912, 0.854347, 0.858385, 0.861996, 0.865003,
+ 0.86646, 0.82184, 0.821897, 0.821674, 0.821592, 0.821429,
+ 0.86842, 0.871631, 0.874676, 0.877554, 0.928498, 0.936229,
+ 0.943903, 0.951517, 0.95907, 0.902802, 0.908617, 0.914903,
+ 0.921194, 0.927466, 0.912617, 0.919099, 0.925592, 0.932094,
+ 0.938605, 0.915914, 0.921739, 0.928803, 0.935927, 0.943095,
+ 0.982139, 0.992066, 1, 1, 0.970056, 0.977633,
+ 0.985279, 0.992996, 1, 0.981505, 0.988024, 0.995008,
+ 1, 1, 0.97652, 0.981778, 0.987072, 0.992403,
+ 0.997772, 0.989569, 0.994141, 0.99874, 1, 1,
+ 0.958503, 0.959695, 0.960888, 0.961952, 0.984313, 0.987439,
+ 0.99058, 0.993734, 0.996902, 0.986424, 0.988754, 0.991091,
+ 0.993435, 0.995786, 0.984205, 0.985709, 0.987216, 0.988726,
+ 0.990238, 0.991754, 0.993272, 0.994792, 0.996316, 0.997843,
+ 0.997771, 0.99948, 1, 1, 0.978729, 0.978557,
+ 0.978385, 0.978213, 0.978042, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 0.984196, 0.983159, 0.982125, 0.981093, 0.980062,
+ 0.991678, 0.991678, 0.991678, 0.991678, 0.991678, 1,
+ 1, 1, 1, 1)"
+          tdata_1to0_min="(1.63161e-011, 2.2246e-011, 2.81759e-011, 3.41058e-011, 4.00356e-011, 4.59655e-011,
+ 5.18954e-011, 5.78253e-011, 6.37551e-011, 6.9685e-011, 7.56149e-011, 8.15448e-011,
+ 8.74746e-011, 9.34045e-011, 9.93344e-011, 1.05264e-010, 1.11194e-010, 1.17124e-010,
+ 1.23054e-010, 1.28984e-010, 1.34914e-010, 1.40843e-010, 1.46773e-010, 1.52703e-010,
+ 1.58633e-010, 1.64563e-010, 1.70493e-010, 1.76423e-010, 1.82353e-010, 1.88282e-010,
+ 1.94212e-010, 2.00142e-010, 2.06072e-010, 2.12002e-010, 2.17932e-010, 2.23862e-010,
+ 2.29792e-010, 2.35721e-010, 2.41651e-010, 2.47581e-010, 2.53511e-010, 2.59441e-010,
+ 2.65371e-010, 2.71301e-010, 2.77231e-010, 2.8316e-010, 2.8909e-010, 2.9502e-010,
+ 3.0095e-010, 3.0688e-010, 3.1281e-010, 3.1874e-010, 3.2467e-010, 3.30599e-010,
+ 3.36529e-010, 3.42459e-010, 3.48389e-010, 3.54319e-010, 3.60249e-010, 3.66179e-010,
+ 3.72109e-010, 3.78038e-010, 3.83968e-010, 3.89898e-010, 3.95828e-010, 4.01758e-010,
+ 4.07688e-010, 4.13618e-010, 4.19548e-010, 4.25477e-010, 4.31407e-010, 4.37337e-010,
+ 4.43267e-010, 4.49197e-010, 4.55127e-010, 4.61057e-010, 4.66987e-010, 4.72916e-010,
+ 4.78846e-010, 4.84776e-010, 4.90706e-010, 4.96636e-010, 5.02566e-010, 5.08496e-010,
+ 5.14426e-010, 5.20355e-010, 5.26285e-010, 5.32215e-010, 5.38145e-010, 5.44075e-010,
+ 5.50005e-010, 5.55935e-010, 5.61865e-010, 5.67794e-010, 5.73724e-010, 5.79654e-010,
+ 5.85584e-010, 5.91514e-010, 5.97444e-010, 6.03374e-010, 6.09304e-010, 6.15233e-010,
+ 6.21163e-010, 6.27093e-010, 6.33023e-010, 6.38953e-010, 6.44883e-010, 6.50813e-010,
+ 6.56743e-010, 6.62672e-010, 6.68602e-010, 6.74532e-010, 6.80462e-010, 6.86392e-010,
+ 6.92322e-010, 6.98252e-010, 7.04182e-010, 7.10111e-010, 7.16041e-010, 7.21971e-010,
+ 7.27901e-010, 7.33831e-010, 7.39761e-010, 7.45691e-010, 7.51621e-010, 7.5755e-010,
+ 7.6348e-010, 7.6941e-010, 7.7534e-010, 7.8127e-010, 7.872e-010, 7.9313e-010,
+ 7.9906e-010, 8.04989e-010, 8.10919e-010, 8.16849e-010, 8.22779e-010, 8.28709e-010,
+ 8.34639e-010, 8.40569e-010, 8.46499e-010, 8.52428e-010, 8.58358e-010, 8.64288e-010,
+ 8.70218e-010, 8.76148e-010, 8.82078e-010, 8.88008e-010, 8.93938e-010, 8.99867e-010,
+ 9.05797e-010, 9.11727e-010, 9.17657e-010, 9.23587e-010, 9.29517e-010, 9.35447e-010,
+ 9.41377e-010, 9.47306e-010, 9.53236e-010, 9.59166e-010, 9.65096e-010, 9.71026e-010,
+ 9.76956e-010, 9.82886e-010, 9.88816e-010, 9.94745e-010, 1.00068e-009, 1.00661e-009,
+ 1.01254e-009, 1.01846e-009, 1.02439e-009, 1.03032e-009, 1.03625e-009, 1.04218e-009,
+ 1.04811e-009, 1.05404e-009, 1.05997e-009, 1.0659e-009, 1.07183e-009, 1.07776e-009,
+ 1.08369e-009, 1.08962e-009, 1.09555e-009, 1.10148e-009, 1.10741e-009, 1.11334e-009,
+ 1.11927e-009, 1.1252e-009, 1.13113e-009, 1.13706e-009, 1.14299e-009, 1.14892e-009,
+ 1.15485e-009, 1.16078e-009, 1.16671e-009, 1.17264e-009, 1.17857e-009, 1.1845e-009,
+ 1.19043e-009, 1.19636e-009, 1.20229e-009, 1.20822e-009)"
+          kdata_1to0_min="(1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 0.944958, 0.941817, 0.939014,
+ 0.936329, 0.933652, 0.928097, 0.926197, 0.924296, 0.922394,
+ 0.920489, 0.918327, 0.916081, 0.742328, 0.734287, 0.726279,
+ 0.718306, 0.710366, 0.5818, 0.572814, 0.563786, 0.554718,
+ 0.545614, 0.432759, 0.422287, 0.411632, 0.400804, 0.390031,
+ 0.357675, 0.345405, 0.33285, 0.319786, 0.306318, 0.299028,
+ 0.281999, 0.263834, 0.245179, 0.224, 0.21373, 0.19043,
+ 0.164822, 0.138767, 0.11283, 0.168453, 0.142421, 0.11653,
+ 0.0898447, 0.064093, 0.12499, 0.101151, 0.0779349, 0.0556811,
+ 0.0329568, 0.116942, 0.0977118, 0.0785584, 0.0587776, 0.0393621,
+ 0.100619, 0.0856291, 0.0698708, 0.0543328, 0.0388455, 0.0738995,
+ 0.0617298, 0.0492707, 0.0366203, 0.0238299, 0.0109021, 0.0561065,
+ 0.0467763, 0.0372812, 0.0274446, 0.0172799, 0.0457196, 0.0381295,
+ 0.0304268, 0.0225745, 0.0145697, 0.0383468, 0.0325389, 0.0266255,
+ 0.0206042, 0.0144643, 0.0365308, 0.0322321, 0.0277894, 0.0232542,
+ 0.0186239, 0.028672, 0.025203, 0.0216809, 0.0181047, 0.0144733,
+ 0.0148853, 0.0116153, 0.00831567, 0.00498609, 0.0016262, 0.0188761,
+ 0.0170186, 0.015139, 0.0132368, 0.0113117, 0.0155086, 0.0140556,
+ 0.0125899, 0.0111111, 0.00961925, 0.0139533, 0.0129102, 0.0118597,
+ 0.0108016, 0.00973602, 0.0114324, 0.0105801, 0.00972376, 0.00886338,
+ 0.00799891, 0.00901914, 0.00830074, 0.00758063, 0.0068588, 0.00613525,
+ 0.00561266, 0.00490209, 0.00419006, 0.00347656, 0.00276158, 0.00173159,
+ 0.000988725, 0.000244458, 0, 0, 0.00391781, 0.00364127,
+ 0.00336415, 0.00308644, 0.00280814, 0.00360153, 0.003408, 0.00321424,
+ 0.00302027, 0.00282607, 0.00282379, 0.00264561, 0.00246717, 0.00228846,
+ 0.00210949, 0.00204093, 0.00187022, 0.00169929, 0.00152814, 0.00135675,
+ 0.00118514, 0.00121595, 0.00106019, 0.000904174, 0.000747895, 0.000591352,
+ 0.00127719, 0.00118284, 0.00108844, 0.000993996, 0.000899505, 0.000727513,
+ 0.000625664, 0.000523821, 0.000421982, 0.000320148, 0.000293503, 0.000198808,
+ 0.000104067, 9.27975e-006, 0, 0.0004531, 0.000407536, 0.000361956,
+ 0.000316359, 0.000270744, 0.000225112, 0)"
+          vdata_min="(-1.8, -1.74, -1.68, -1.62, -1.56, -1.5,
+ -1.44, -1.38, -1.32, -1.26, -1.2, -1.14,
+ -1.08, -1.02, -0.96, -0.9, -0.84, -0.78,
+ -0.72, -0.66, -0.6, -0.54, -0.48, -0.42,
+ -0.36, -0.3, -0.24, -0.18, -0.12, -0.06,
+ 0, 0.06, 0.12, 0.18, 0.24, 0.3,
+ 0.36, 0.42, 0.48, 0.54, 0.6, 0.66,
+ 0.72, 0.78, 0.84, 0.9, 0.96, 1.02,
+ 1.08, 1.14, 1.2, 1.26, 1.32, 1.38,
+ 1.44, 1.5, 1.56, 1.62, 1.68, 1.74,
+ 1.8, 1.86, 1.92, 1.98, 2.04, 2.1,
+ 2.16, 2.22, 2.28, 2.34, 2.4, 2.46,
+ 2.52, 2.58, 2.64, 2.7, 2.76, 2.82,
+ 2.88, 2.94, 3, 3.06, 3.12, 3.18,
+ 3.24, 3.3, 3.36, 3.42, 3.48, 3.54,
+ 3.6)"
+          idata_min="(-2.394, -2.235, -2.075, -1.915, -1.756, -1.596,
+ -1.437, -1.277, -1.118, -0.9586, -0.7993, -0.6403,
+ -0.4841, -0.3375, -0.2096, -0.1333, -0.1135, -0.1032,
+ -0.09427, -0.08574, -0.07761, -0.06996, -0.06286, -0.05631,
+ -0.05017, -0.04422, -0.03837, -0.03258, -0.02687, -0.02127,
+ -0.01578, -0.01053, -0.005574, -0.0009032, 0.003482, 0.007583,
+ 0.0114, 0.01494, 0.0182, 0.02119, 0.0239, 0.02632,
+ 0.02844, 0.03027, 0.03189, 0.03338, 0.03481, 0.0362,
+ 0.03759, 0.03898, 0.04039, 0.04181, 0.04324, 0.0447,
+ 0.04617, 0.04766, 0.04918, 0.05073, 0.0523, 0.0539,
+ 0.05554, 0.05721, 0.05887, 0.06051, 0.06215, 0.06379,
+ 0.06553, 0.06774, 0.07132, 0.07727, 0.08581, 0.09653,
+ 0.109, 0.1233, 0.143, 0.1988, 0.4466, 0.8356,
+ 1.244, 1.664, 2.088, 2.513, 2.938, 3.364,
+ 3.79, 4.216, 4.641, 5.067, 5.493, 5.919,
+ 6.346)"
+          tdata_0to1_max="(7.19709e-011, 7.82209e-011, 8.44709e-011, 9.07209e-011, 9.69709e-011, 1.03221e-010,
+ 1.09471e-010, 1.15721e-010, 1.21971e-010, 1.28221e-010, 1.34471e-010, 1.40721e-010,
+ 1.46971e-010, 1.53221e-010, 1.59471e-010, 1.65721e-010, 1.71971e-010, 1.78221e-010,
+ 1.84471e-010, 1.90721e-010, 1.96971e-010, 2.03221e-010, 2.09471e-010, 2.15721e-010,
+ 2.21971e-010, 2.28221e-010, 2.34471e-010, 2.40721e-010, 2.46971e-010, 2.53221e-010,
+ 2.59471e-010, 2.65721e-010, 2.71971e-010, 2.78221e-010, 2.84471e-010, 2.90721e-010,
+ 2.96971e-010, 3.03221e-010, 3.09471e-010, 3.15721e-010, 3.21971e-010, 3.28221e-010,
+ 3.34471e-010, 3.40721e-010, 3.46971e-010, 3.53221e-010, 3.59471e-010, 3.65721e-010,
+ 3.71971e-010, 3.78221e-010, 3.84471e-010, 3.90721e-010, 3.96971e-010, 4.03221e-010,
+ 4.09471e-010, 4.15721e-010, 4.21971e-010, 4.28221e-010, 4.34471e-010, 4.40721e-010,
+ 4.46971e-010, 4.53221e-010, 4.59471e-010, 4.65721e-010, 4.71971e-010, 4.78221e-010,
+ 4.84471e-010, 4.90721e-010, 4.96971e-010, 5.03221e-010, 5.09471e-010, 5.15721e-010,
+ 5.21971e-010, 5.28221e-010, 5.34471e-010, 5.40721e-010, 5.46971e-010, 5.53221e-010,
+ 5.59471e-010, 5.65721e-010, 5.71971e-010, 5.78221e-010, 5.84471e-010, 5.90721e-010,
+ 5.96971e-010, 6.03221e-010, 6.09471e-010, 6.15721e-010, 6.21971e-010, 6.28221e-010,
+ 6.34471e-010, 6.40721e-010, 6.46971e-010, 6.53221e-010, 6.59471e-010, 6.65721e-010,
+ 6.71971e-010, 6.78221e-010, 6.84471e-010, 6.90721e-010, 6.96971e-010, 7.03221e-010,
+ 7.09471e-010, 7.15721e-010, 7.21971e-010, 7.28221e-010, 7.34471e-010, 7.40721e-010,
+ 7.46971e-010, 7.53221e-010, 7.59471e-010, 7.65721e-010, 7.71971e-010, 7.78221e-010,
+ 7.84471e-010, 7.90721e-010, 7.96971e-010, 8.03221e-010, 8.09471e-010, 8.15721e-010,
+ 8.21971e-010, 8.28221e-010, 8.34471e-010, 8.40721e-010, 8.46971e-010, 8.53221e-010,
+ 8.59471e-010, 8.65721e-010, 8.71971e-010, 8.78221e-010, 8.84471e-010, 8.90721e-010,
+ 8.96971e-010, 9.03221e-010, 9.09471e-010, 9.15721e-010, 9.21971e-010, 9.28221e-010,
+ 9.34471e-010, 9.40721e-010, 9.46971e-010, 9.53221e-010, 9.59471e-010, 9.65721e-010,
+ 9.71971e-010, 9.78221e-010, 9.84471e-010, 9.90721e-010, 9.96971e-010, 1.00322e-009,
+ 1.00947e-009, 1.01572e-009, 1.02197e-009, 1.02822e-009, 1.03447e-009, 1.04072e-009,
+ 1.04697e-009, 1.05322e-009, 1.05947e-009, 1.06572e-009, 1.07197e-009, 1.07822e-009,
+ 1.08447e-009, 1.09072e-009, 1.09697e-009, 1.10322e-009, 1.10947e-009, 1.11572e-009,
+ 1.12197e-009, 1.12822e-009, 1.13447e-009, 1.14072e-009, 1.14697e-009, 1.15322e-009,
+ 1.15947e-009, 1.16572e-009, 1.17197e-009, 1.17822e-009, 1.18447e-009, 1.19072e-009,
+ 1.19697e-009, 1.20322e-009, 1.20947e-009, 1.21572e-009, 1.22197e-009, 1.22822e-009,
+ 1.23447e-009, 1.24072e-009, 1.24697e-009, 1.25322e-009, 1.25947e-009, 1.26572e-009,
+ 1.27197e-009, 1.27822e-009, 1.28447e-009, 1.29072e-009, 1.29697e-009, 1.30322e-009,
+ 1.30947e-009, 1.31572e-009, 1.32197e-009, 1.32822e-009)"
+          kdata_0to1_max="(0, 0.00144844, 0.00161591, 0.00178283, 0.00194921, 0.00211506,
+ 0.0087038, 0.00937234, 0.0100361, 0.0106951, 0.0113493, 0.0221732,
+ 0.0235462, 0.0248913, 0.0262091, 0.027512, 0.0384896, 0.040387,
+ 0.0422566, 0.0440992, 0.0459152, 0.0477052, 0.0909226, 0.0947716,
+ 0.0985008, 0.102115, 0.10562, 0.151672, 0.156561, 0.161263,
+ 0.165788, 0.170143, 0.231451, 0.237879, 0.244041, 0.249991,
+ 0.255738, 0.306646, 0.314487, 0.322133, 0.329544, 0.346723,
+ 0.354268, 0.361647, 0.368849, 0.375871, 0.436727, 0.446473,
+ 0.456075, 0.465528, 0.47489, 0.508024, 0.518296, 0.528421,
+ 0.538431, 0.548284, 0.578952, 0.589365, 0.599555, 0.609511,
+ 0.619187, 0.661993, 0.673295, 0.684356, 0.695153, 0.695174,
+ 0.703634, 0.711667, 0.719248, 0.725866, 0.705895, 0.708557,
+ 0.710598, 0.711564, 0.710588, 0.813801, 0.819259, 0.824199,
+ 0.827163, 0.82912, 0.854347, 0.858385, 0.861996, 0.865003,
+ 0.86646, 0.82184, 0.821897, 0.821674, 0.821592, 0.821429,
+ 0.86842, 0.871631, 0.874676, 0.877554, 0.928498, 0.936229,
+ 0.943903, 0.951517, 0.95907, 0.902802, 0.908617, 0.914903,
+ 0.921194, 0.927466, 0.912617, 0.919099, 0.925592, 0.932094,
+ 0.938605, 0.915914, 0.921739, 0.928803, 0.935927, 0.943095,
+ 0.982139, 0.992066, 1, 1, 0.970056, 0.977633,
+ 0.985279, 0.992996, 1, 0.981505, 0.988024, 0.995008,
+ 1, 1, 0.97652, 0.981778, 0.987072, 0.992403,
+ 0.997772, 0.989569, 0.994141, 0.99874, 1, 1,
+ 0.958503, 0.959695, 0.960888, 0.961952, 0.984313, 0.987439,
+ 0.99058, 0.993734, 0.996902, 0.986424, 0.988754, 0.991091,
+ 0.993435, 0.995786, 0.984205, 0.985709, 0.987216, 0.988726,
+ 0.990238, 0.991754, 0.993272, 0.994792, 0.996316, 0.997843,
+ 0.997771, 0.99948, 1, 1, 0.978729, 0.978557,
+ 0.978385, 0.978213, 0.978042, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 0.984196, 0.983159, 0.982125, 0.981093, 0.980062,
+ 0.991678, 0.991678, 0.991678, 0.991678, 0.991678, 1,
+ 1, 1, 1, 1)"
+          tdata_1to0_max="(1.63161e-011, 2.2246e-011, 2.81759e-011, 3.41058e-011, 4.00356e-011, 4.59655e-011,
+ 5.18954e-011, 5.78253e-011, 6.37551e-011, 6.9685e-011, 7.56149e-011, 8.15448e-011,
+ 8.74746e-011, 9.34045e-011, 9.93344e-011, 1.05264e-010, 1.11194e-010, 1.17124e-010,
+ 1.23054e-010, 1.28984e-010, 1.34914e-010, 1.40843e-010, 1.46773e-010, 1.52703e-010,
+ 1.58633e-010, 1.64563e-010, 1.70493e-010, 1.76423e-010, 1.82353e-010, 1.88282e-010,
+ 1.94212e-010, 2.00142e-010, 2.06072e-010, 2.12002e-010, 2.17932e-010, 2.23862e-010,
+ 2.29792e-010, 2.35721e-010, 2.41651e-010, 2.47581e-010, 2.53511e-010, 2.59441e-010,
+ 2.65371e-010, 2.71301e-010, 2.77231e-010, 2.8316e-010, 2.8909e-010, 2.9502e-010,
+ 3.0095e-010, 3.0688e-010, 3.1281e-010, 3.1874e-010, 3.2467e-010, 3.30599e-010,
+ 3.36529e-010, 3.42459e-010, 3.48389e-010, 3.54319e-010, 3.60249e-010, 3.66179e-010,
+ 3.72109e-010, 3.78038e-010, 3.83968e-010, 3.89898e-010, 3.95828e-010, 4.01758e-010,
+ 4.07688e-010, 4.13618e-010, 4.19548e-010, 4.25477e-010, 4.31407e-010, 4.37337e-010,
+ 4.43267e-010, 4.49197e-010, 4.55127e-010, 4.61057e-010, 4.66987e-010, 4.72916e-010,
+ 4.78846e-010, 4.84776e-010, 4.90706e-010, 4.96636e-010, 5.02566e-010, 5.08496e-010,
+ 5.14426e-010, 5.20355e-010, 5.26285e-010, 5.32215e-010, 5.38145e-010, 5.44075e-010,
+ 5.50005e-010, 5.55935e-010, 5.61865e-010, 5.67794e-010, 5.73724e-010, 5.79654e-010,
+ 5.85584e-010, 5.91514e-010, 5.97444e-010, 6.03374e-010, 6.09304e-010, 6.15233e-010,
+ 6.21163e-010, 6.27093e-010, 6.33023e-010, 6.38953e-010, 6.44883e-010, 6.50813e-010,
+ 6.56743e-010, 6.62672e-010, 6.68602e-010, 6.74532e-010, 6.80462e-010, 6.86392e-010,
+ 6.92322e-010, 6.98252e-010, 7.04182e-010, 7.10111e-010, 7.16041e-010, 7.21971e-010,
+ 7.27901e-010, 7.33831e-010, 7.39761e-010, 7.45691e-010, 7.51621e-010, 7.5755e-010,
+ 7.6348e-010, 7.6941e-010, 7.7534e-010, 7.8127e-010, 7.872e-010, 7.9313e-010,
+ 7.9906e-010, 8.04989e-010, 8.10919e-010, 8.16849e-010, 8.22779e-010, 8.28709e-010,
+ 8.34639e-010, 8.40569e-010, 8.46499e-010, 8.52428e-010, 8.58358e-010, 8.64288e-010,
+ 8.70218e-010, 8.76148e-010, 8.82078e-010, 8.88008e-010, 8.93938e-010, 8.99867e-010,
+ 9.05797e-010, 9.11727e-010, 9.17657e-010, 9.23587e-010, 9.29517e-010, 9.35447e-010,
+ 9.41377e-010, 9.47306e-010, 9.53236e-010, 9.59166e-010, 9.65096e-010, 9.71026e-010,
+ 9.76956e-010, 9.82886e-010, 9.88816e-010, 9.94745e-010, 1.00068e-009, 1.00661e-009,
+ 1.01254e-009, 1.01846e-009, 1.02439e-009, 1.03032e-009, 1.03625e-009, 1.04218e-009,
+ 1.04811e-009, 1.05404e-009, 1.05997e-009, 1.0659e-009, 1.07183e-009, 1.07776e-009,
+ 1.08369e-009, 1.08962e-009, 1.09555e-009, 1.10148e-009, 1.10741e-009, 1.11334e-009,
+ 1.11927e-009, 1.1252e-009, 1.13113e-009, 1.13706e-009, 1.14299e-009, 1.14892e-009,
+ 1.15485e-009, 1.16078e-009, 1.16671e-009, 1.17264e-009, 1.17857e-009, 1.1845e-009,
+ 1.19043e-009, 1.19636e-009, 1.20229e-009, 1.20822e-009)"
+          kdata_1to0_max="(1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 1, 1, 1,
+ 1, 1, 1, 0.944958, 0.941817, 0.939014,
+ 0.936329, 0.933652, 0.928097, 0.926197, 0.924296, 0.922394,
+ 0.920489, 0.918327, 0.916081, 0.742328, 0.734287, 0.726279,
+ 0.718306, 0.710366, 0.5818, 0.572814, 0.563786, 0.554718,
+ 0.545614, 0.432759, 0.422287, 0.411632, 0.400804, 0.390031,
+ 0.357675, 0.345405, 0.33285, 0.319786, 0.306318, 0.299028,
+ 0.281999, 0.263834, 0.245179, 0.224, 0.21373, 0.19043,
+ 0.164822, 0.138767, 0.11283, 0.168453, 0.142421, 0.11653,
+ 0.0898447, 0.064093, 0.12499, 0.101151, 0.0779349, 0.0556811,
+ 0.0329568, 0.116942, 0.0977118, 0.0785584, 0.0587776, 0.0393621,
+ 0.100619, 0.0856291, 0.0698708, 0.0543328, 0.0388455, 0.0738995,
+ 0.0617298, 0.0492707, 0.0366203, 0.0238299, 0.0109021, 0.0561065,
+ 0.0467763, 0.0372812, 0.0274446, 0.0172799, 0.0457196, 0.0381295,
+ 0.0304268, 0.0225745, 0.0145697, 0.0383468, 0.0325389, 0.0266255,
+ 0.0206042, 0.0144643, 0.0365308, 0.0322321, 0.0277894, 0.0232542,
+ 0.0186239, 0.028672, 0.025203, 0.0216809, 0.0181047, 0.0144733,
+ 0.0148853, 0.0116153, 0.00831567, 0.00498609, 0.0016262, 0.0188761,
+ 0.0170186, 0.015139, 0.0132368, 0.0113117, 0.0155086, 0.0140556,
+ 0.0125899, 0.0111111, 0.00961925, 0.0139533, 0.0129102, 0.0118597,
+ 0.0108016, 0.00973602, 0.0114324, 0.0105801, 0.00972376, 0.00886338,
+ 0.00799891, 0.00901914, 0.00830074, 0.00758063, 0.0068588, 0.00613525,
+ 0.00561266, 0.00490209, 0.00419006, 0.00347656, 0.00276158, 0.00173159,
+ 0.000988725, 0.000244458, 0, 0, 0.00391781, 0.00364127,
+ 0.00336415, 0.00308644, 0.00280814, 0.00360153, 0.003408, 0.00321424,
+ 0.00302027, 0.00282607, 0.00282379, 0.00264561, 0.00246717, 0.00228846,
+ 0.00210949, 0.00204093, 0.00187022, 0.00169929, 0.00152814, 0.00135675,
+ 0.00118514, 0.00121595, 0.00106019, 0.000904174, 0.000747895, 0.000591352,
+ 0.00127719, 0.00118284, 0.00108844, 0.000993996, 0.000899505, 0.000727513,
+ 0.000625664, 0.000523821, 0.000421982, 0.000320148, 0.000293503, 0.000198808,
+ 0.000104067, 9.27975e-006, 0, 0.0004531, 0.000407536, 0.000361956,
+ 0.000316359, 0.000270744, 0.000225112, 0)"
+          vdata_max="(-1.8, -1.74, -1.68, -1.62, -1.56, -1.5,
+ -1.44, -1.38, -1.32, -1.26, -1.2, -1.14,
+ -1.08, -1.02, -0.96, -0.9, -0.84, -0.78,
+ -0.72, -0.66, -0.6, -0.54, -0.48, -0.42,
+ -0.36, -0.3, -0.24, -0.18, -0.12, -0.06,
+ 0, 0.06, 0.12, 0.18, 0.24, 0.3,
+ 0.36, 0.42, 0.48, 0.54, 0.6, 0.66,
+ 0.72, 0.78, 0.84, 0.9, 0.96, 1.02,
+ 1.08, 1.14, 1.2, 1.26, 1.32, 1.38,
+ 1.44, 1.5, 1.56, 1.62, 1.68, 1.74,
+ 1.8, 1.86, 1.92, 1.98, 2.04, 2.1,
+ 2.16, 2.22, 2.28, 2.34, 2.4, 2.46,
+ 2.52, 2.58, 2.64, 2.7, 2.76, 2.82,
+ 2.88, 2.94, 3, 3.06, 3.12, 3.18,
+ 3.24, 3.3, 3.36, 3.42, 3.48, 3.54,
+ 3.6)"
+          idata_max="(-2.394, -2.235, -2.075, -1.915, -1.756, -1.596,
+ -1.437, -1.277, -1.118, -0.9586, -0.7993, -0.6403,
+ -0.4841, -0.3375, -0.2096, -0.1333, -0.1135, -0.1032,
+ -0.09427, -0.08574, -0.07761, -0.06996, -0.06286, -0.05631,
+ -0.05017, -0.04422, -0.03837, -0.03258, -0.02687, -0.02127,
+ -0.01578, -0.01053, -0.005574, -0.0009032, 0.003482, 0.007583,
+ 0.0114, 0.01494, 0.0182, 0.02119, 0.0239, 0.02632,
+ 0.02844, 0.03027, 0.03189, 0.03338, 0.03481, 0.0362,
+ 0.03759, 0.03898, 0.04039, 0.04181, 0.04324, 0.0447,
+ 0.04617, 0.04766, 0.04918, 0.05073, 0.0523, 0.0539,
+ 0.05554, 0.05721, 0.05887, 0.06051, 0.06215, 0.06379,
+ 0.06553, 0.06774, 0.07132, 0.07727, 0.08581, 0.09653,
+ 0.109, 0.1233, 0.143, 0.1988, 0.4466, 0.8356,
+ 1.244, 1.664, 2.088, 2.513, 2.938, 3.364,
+ 3.79, 4.216, 4.641, 5.067, 5.493, 5.919,
+ 6.346)"
+ PORT: a_signal
+       a_PuRef
+       d_pullup_control

.model ibis_ktiv(icx_behavioral) MACRO LANG=VHDLAMS LIB=icxbase
.ends MODEL_U3_1

