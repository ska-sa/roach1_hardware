* OrCAD Model Editor - Version 10.1
*
*  AD8027devel Spice Macro-model           ADI
*John Ardizzoni 
*8027_3/3/04
*  Copyright 2004 by Analog Devices, Inc.
*
* Refer to "README.DOC" file for License Statement.
* Use of this model indicates your acceptance with
* the terms and provisions in the License Statement.
*
* The following parameters are accurately modeled;
*
*    open loop gain and phase vs frequency
*    output clamping voltage and current
*    input common mode range
*    CMRR vs freq
*    I bias vs Vcm in    
*    Slew rate
*    Output currents are reflected to V supplies
*
*    Vos is static and will not vary with Vcm in
*    Step response is modeled at unity gain w/1k load 
*
*    Distortion and noise are not characterized
*
*    Node assignments
*                non-inverting input
*                | inverting input
*                | | positive supply
*                | | |  negative supply
*                | | |  |  output
*                | | |  |  |
.SUBCKT AD8027  1 2 99 50 61   

***** Input bias current source

ecm 20 0 3 97 1 
d1 20 21 dx
d2 23 20 dx
v3 21 22 -0.9
v4 24 23 -0.9
r20 22 0 100
r21 24 0 100
f1 0 25 v3 1 
f2 25 0 v4 1
r22 25 0 1k
d3 25 26 dx
d4 27 25 dx
v5 26 0 .2
v6 0 27 .2
g1 1 0 25 0 3.8e-6
g2 2 0 25 0 3.8e-6

***** Input Stage

R1 1 3 3Meg
R2 3 2 3Meg
C1 1 2 2pf
R3 1 98 40e6
R4 2 98 40e6 
r9 15 7 29.45
r10 16 7 29.45
q1 5 1 15 qn1
q2 6 4 16 qn1
r5 99 5 81.45
r6 99 6 81.45
cp 5 6 4pf
ib3 7 50 1e-3
eos 2 4 poly(1) (1501,98) 0.24e-3 1 
*Vos 2 4 .24e-3

***** dummy first stage (pnp) for correct bias current

ib4 81 99 1e-3
r11 82 81 1015
r12 83 81 1015
q3 84 1 82 qp1 
q4 85 4 83 qp1
r13 50 84 1515
r14 50 85 1515

***** gain stage/pole at 1000hz/clamp circuitry

g3 99 31 6 5 .012
g4 31 50 5 6 .012
r7 99 31 15.915e6
r8 31 50 15.915e6
c3 99 31 10e-12
c4 31 50 10e-12
vc1 99 45 -0.85
vc2 46 50 -0.85
dc1 31 45 dx
dc2 46 31 dx

***** pole/zero 6KHz/8KHz

g100 99 42 31 98 1u
g101 42 50 98 31 1u
r300 99 42 1e6
r301 42 50 1e6
R3000 99 3000 3E6
R3001 50 3001 3E6
C1000 3000 42 19.89e-12
C1001 42 3001 19.89e-12

****zero/pole 112MHz/300M
g51 99 331 42 0 1u
g61 331 50 0 42 1u
Rg11 99 341 1.68e6
Rg21 341 331 1e6
Lg11 99 341 .89e-3 
Rg31 351 331 1e6
Rg41 351 50 1.68e6
Lg21 351 50 .89e-3

***** internal reference
rdiv1 99 97 100k
rdiv2 97 50 100k
Eref 98 0 97 0 1
rref 98 0 1e6

****Common mode gain and 10KHz zero network
gcm1 99 105 3 98 2.4e-12
gcm2 105 50 98 3 2.4e-12
l1cm 99 103 10.5
l2cm 106 50 10.5
racm1 103 105 1e6
racm2 105 106 1e6

*****Common Mode gain Zero at 16MHz
gcmz1 99 145 105 98 1u
gcmz2 145 50 98 105 1u
lcmz1 99 140 9.94e-3
lcmz2 141 50 9.94e-3
racmz1 140 145 1e6
racmz2 145 141 1e6

***** Common Mode Gain Pole at 70MHz 

gccm1 99 150 145 98 1u
gccm2 150 50 98 145 1u
rcmpole1 99 150 1e6
rcmpole2 150 50 1e6
cmpole1 99 150 2.27e-15
cmpole2 150 50 2.27e-15

***** Common Mode Pole at 150MHz 

gccm11 99 1501 150 98 1u
gccm21 150 50 98 150 1u
rcmpole11 99 1501 1e6
rcmpole21 1501 50 1e6
cmpole11 99 1501 1.06e-15
cmpole21 1501 50 1.06e-15

***** buffer to output stage

gbuf 98 32 331 98 1e-4
re1 32 98 10k

***** output stage

fo1 98 110 vcd 1
do1 110 111 dx
do2 112 110 dx
vi1 111 98 0
vi2 98 112 0

fsy 99 50 poly(2) vi1 vi2 6.0e-3 1 1

go3 60 99 99 32 50
go4 50 60 32 50 50
r03 60 99 .02
r04 60 50 .02
vcd 60 62 0
lo1 62 61 .01u
*ro1 62 61 .01
ro2 61 98 1e9
do5 32 70 dx
do6 71 32 dx
vo1 70 60 -0.699
vo2 60 71 -0.699

.model dx d(is=1e-15)
.model qn1 npn(bf=91 vaf=100)
.model qp1 pnp(bf=2500 vaf=60)
.ends


