* OP176G SPICE Macro-model             11/93, Rev. A
*                                       ARG / PMI
*
* This version of the OP-176 model simulates the worst-case
* parameters of the 'G' grade.  The worst-case parameters
* used correspond to those in the data sheet.
*
* Copyright 1992 by Analog Devices
*
* Refer to "README.DOC" file for License Statement.  Use of this model
* indicates your acceptance with the terms and provisions in the License
* Statement.
*
* Node assignments
*               non-inverting input
*               | inverting input
*               | | positive supply
*               | | |  negative supply
*               | | |  |  output
*               | | |  |  |
*               | | |  |  |
.SUBCKT OP176G  1 2 99 50 34
*
* INPUT STAGE & POLE AT 100MHZ
*
R3   5 51     1.492
R4   6 51     1.492
CIN  1  2     3.7E-12
CM1  1 98     7.5E-12
CM2  2 98     7.5E-12
C2   5  6     320E-12
I1   97 4     100E-3
IOS  1  2     25E-9
EOS  9  3     POLY(1)  (26,28)  1E-3  1
Q1   5  2  7  QX
Q2   6  9  8  QX
R5   7  4     0.975
R6   8  4     0.975
D1   2 36     DZ
D2   1 36     DZ
EN   3  1     (10,0)  1
GN1  0  2     (13,0)  1E-3
GN2  0  1     (16,0)  1E-3
*
EREF 98 0     (28,0)  1
EP   97 0     (99,0)  1
EM   51 0     (50,0)  1
*
* VOLTAGE NOISE SOURCE
*
DN1  35 10    DEN
DN2  10 11    DEN
VN1  35  0    DC 2
VN2  0  11    DC 2
*
* CURRENT NOISE SOURCE
*
DN3  12 13    DIN
DN4  13 14    DIN
VN3  12  0    DC 2
VN4  0  14    DC 2
*
* CURRENT NOISE SOURCE
*
DN5  15 16    DIN
DN6  16 17    DIN
VN5  15  0    DC 2
VN6  0  17    DC 2
*
* GAIN STAGE & DOMINANT POLE AT 64HZ
*
R7  18 98     373.019E3
C3  18 98     6.667E-9
G1  98 18     (5,6)  670.206E-3
V2  97 19     1.82
V3  20 51     1.82
D3  18 19     DX
D4  20 18     DX
*
* POLE/ZERO PAIR AT 1.5MHZ/2.7MHZ
*
R8  21 98     1E3
R9  21 22     1.25E3
C4  22 98     47.2E-12
G2  98 21     (18,28)  1E-3
*
* POLE AT 100MHZ
*
R10 23 98     1
C5  23 98     1.59E-9
G3  98 23     (21,28)  1
*
* POLE AT 100MHZ
*
R11 24 98     1
C6  24 98     1.59E-9
G4  98 24     (23,28)  1
*
* COMMON-MODE GAIN NETWORK WITH ZERO AT 20KHZ
*
R12 25 26     1E6
C7  25 26     3.183E-12
R13 26 98     1
E2  25 98     POLY(2) (1,98) (2,98) 0 50 50
*
* POLE AT 100MHZ
*
R14 27 98     1
C8  27 98     1.59E-9
G5  98 27     (24,28)  1
*
* OUTPUT STAGE
*
R15 28 99     28E3
R16 28 50     28E3
C9  28 50     1E-6
ISY 99 50     1.964E-3
R17 29 99     100
R18 29 50     100
L2  29 34     1E-9
G6  32 50     (27,29)  10E-3
G7  33 50     (29,27)  10E-3
G8  29 99     (99,27)  10E-3
G9  50 29     (27,50)  10E-3
V4  30 29     0.475
V5  29 31     0.475
F1  29  0     V4  1
F2  0  29     V5  1
D5  27 30     DX
D6  31 27     DX
D7  99 32     DX
D8  99 33     DX
D9  50 32     DY
D10 50 33     DY
*
* MODELS USED
*
.MODEL QX PNP(BF=142.857E3)
.MODEL DX   D(IS=1E-12)
.MODEL DY   D(IS=1E-15 BV=50)
.MODEL DZ   D(IS=1E-15 BV=7.0)
.MODEL DEN  D(IS=1E-12 RS=4.35K KF=1.95E-15 AF=1)
.MODEL DIN  D(IS=1E-12 RS=268 KF=1.08E-15 AF=1)
.ENDS
