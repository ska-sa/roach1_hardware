* BUF04 SPICE Macro-model                  7/93, Rev. A   
*                                           JCB / PMI
*
* Copyright 1993 by Analog Devices, Inc.
*
* Refer to "README.DOC" file for License Statement.
* Use of this model indicates your acceptance with
* the terms and provisions in the License Statement.
*
* Node assignments
*                non-inverting input
*                | positive supply
*                | |  negative supply
*                | |  |  output
*                | |  |  |
*                | |  |  |
.SUBCKT BUF04    1 99 50 6
*
* INPUT STAGE
*
R1   99  8     200
R2   10 50     200
V1   99  9     4.4
D1   9   8     DX
V2   11 50     4.4
D2   10 11     DX
I1   99  5     1.8E-3
I2   4  50     1.8E-3
Q1   50  3  5  QP
Q2   99  3  4  QN
Q3   8  61 30  QN
Q4   10  7 30  QP
R3   5  61     50E3
R4   4   7     50E3
CP1  61 99     14E-15
CP2  7  50     14E-15
RFB  6   2     100
*
* INPUT ERROR SOURCES
* 
IB1  99  1     0.7E-6
VOS  3   1     0.3E-3
LS1  30  2     1E-9
CS1  99  2     2.0E-12
CS2  99  1     3.0E-12
*
EREF 97  0     22  0  1
*
* TRANSCONDUCTANCE STAGE
*
R5   12 97     365E3
C3   12 97     8E-12
G1   97 12     99  8  5E-3
G2   12 97     10 50  5E-3
E3   13 97     POLY(1) 99 97  -2.5  1.1 
E4   97 14     POLY(1) 97 50  -2.5  1.1
D3   12 13     DX
D4   14 12     DX
R6   12 15     200
C2   15  6     20E-12
*
* POLE AT 200 MHZ
*
R11 20 97     1E6
C7  20 97     0.759E-15
G7  97 20     12 22  1E-6
*
* POLE AT 200 MHZ
*
R12 21 97     1E6
C8  21 97     0.759E-15
G8  97 21     20 22  1E-6
*
* OUTPUT STAGE
*
FSY 99 50     POLY(2) V7 V8 1.85E-3 1 1
R13 22 99     16.67E3
R14 22 50     16.67E3
R15 27 99     80
R16 27 50     80
L2  27  6     10E-9
G11 27 99     99 21  12.5E-3
G12 50 27     21 50  12.5E-3
V5  23 27     3.3
V6  27 24     3.3
D5  21 23     DX
D6  24 21     DX
G10 97 70     27 21 12.5E-3
D7  70 71     DX
D8  72 70     DX
V7  71 97     DC 0
V8  97 72     DC 0
*
* MODELS USED
*
.MODEL QN   NPN(BF=1000 IS=1E-15)
.MODEL QP   PNP(BF=1000 IS=1E-15)
.MODEL DX   D(IS=1E-15)
.ENDS
