* AD8591/92/94 SPICE Macro-model Typical Values
* 6/98, Ver. 1
* TAM / ADSC
*
* Copyright 1998 by Analog Devices
*
* Refer to "README.DOC" file for License Statement.  Use of this
* model indicates your acceptance of the terms and provisions in
* the License Statement.
*
* Node Assignments
*		noninverting input
*		|	inverting input
*		|	|	 positive supply
*		|	|	 |	 negative supply
*		|	|	 |	 |	 output
*		|	|	 |	 |	 |	shutdown
*		|	|	 |	 |	 |	|
.SUBCKT AD8592	1	2	99	50	45	80
*
* INPUT STAGE
*
M1   4  1 3 3 PIX L=0.8E-6 W=125E-6
M2   6  7 3 3 PIX L=0.8E-6 W=125E-6
RC1  4 50 4E3
RC2  6 50 4E3
C1   4  6 2E-12
I1  99  8 100E-6

M3  10  1 12 12 NIX L=0.8E-6 W=125E-6
M4  11  7 12 12 NIX L=0.8E-6 W=125E-6
RC3 10 99 4E3
RC4 11 99 4E3
C2  10 11 2E-12
I2  13 50 100E-6

EOS  7  2 POLY(3) (21,98) (73,98) (61,0) 1E-3 0 0 1
IOS  1  2 2.5E-12
V1  99  9 0.9
D1   3  9 DX
V2  14 50 0.9
D2  14 12 DX
S1   3  8 (82,98) SOPEN
S2  99  8 (98,82) SCLOSE
S3  12 13 (82,98) SOPEN
S4  13 50 (98,82) SCLOSE
*
* CMRR 64dB, ZERO AT 20kHz
*
ECM1 20 98 POLY(2) (1,98) (2,98) 0 .5 .5
RCM1 20 21 79.6E3
CCM1 20 21 100E-12
RCM2 21 98 50
*
* PSRR=80dB, ZERO AT 200Hz
*
RPS1 70  0 1E6
RPS2 71  0 1E6
CPS1 99 70 1E-5
CPS2 50 71 1E-5
EPSY 98 72 POLY(2) (70,0) (0,71) 0 1 1
RPS3 72 73 1.59E6
CPS3 72 73 500E-12
RPS4 73 98 80
*
* INTERNAL VOLTAGE REFERENCE
*
EREF 98  0 POLY(2) (99,0) (50,0) 0 .5 .5
GSY  99 50 POLY(1) (99,50) 20E-6 10E-7
*
* SHUTDOWN SECTION
*
E1 81 98 (80,50) 1
R1 81 82 1E3
C3 82 98 1E-9
*
* VOLTAGE NOISE REFERENCE OF 30nV/rt(Hz)
*
VN1 60 0 0
RN1 60 0 16.45E-3
HN  61 0 VN1 30
RN2 61 0 1
*
* GAIN STAGE
*
G2  98 30 POLY(2) (4,6) (10,11) 0 2.19E-5 2.19E-5
R2  30 98 13E6
CF  45 30 5E-12
S5  30 98 (98,82) SCLOSE
D3  30 31 DX
D4  32 30 DX
V3  99 31 0.6
V4  32 50 0.6
*
* OUTPUT STAGE
*
M5  45 46 99 99 POX L=0.8E-6 W=16E-3
M6  45 47 50 50 NOX L=0.8E-6 W=16E-3
EG1 99 48 POLY(1) (98,30) 1.06 1
EG2 49 50 POLY(1) (30,98) 1.05 1
RG1 48 46 10E3
RG2 49 47 10E3
S6  46 99 (98,82) SCLOSE
S7  47 50 (98,82) SCLOSE
*
* MODELS
*
.MODEL PIX PMOS (LEVEL=2,KP=20E-6,VTO=-0.7,LAMBDA=0.01,KF=1E-31)
.MODEL NIX NMOS (LEVEL=2,KP=20E-6,VTO=0.7,LAMBDA=0.01,KF=1E-31)
.MODEL POX PMOS (LEVEL=2,KP=8E-6,VTO=-1,LAMBDA=0.067)
.MODEL NOX NMOS (LEVEL=2,KP=13.4E-6,VTO=1,LAMBDA=0.067)
.MODEL SOPEN VSWITCH(VON=2.4,VOFF=0.8,RON=10,ROFF=1E9)
.MODEL SCLOSE VSWITCH(VON=-0.8,VOFF=-2.4,RON=10,ROFF=1E9)
.MODEL DX D(IS=1E-14)
.ENDS AD8592