* ADG407B SPICE Macro-model                10/95, Rev. D
*                                           WF / ADSC
*
* Revision History: NONE
*
*       NOTE: This model was setup with Maximum leakage currents
*               at +85C for ADG407B
* Copyright 1995 by Analog Devices, Inc.
*
* Refer to "README.DOC" file for License Statement.  Use of this 
* model indicates your acceptance with the terms and provisions 
* in the License Statement.
*
* Node assignments
* 19 - S1A, 20 - S2A, 21 - S3A, 22 - S4A, 23 - S5A, 24 - S6A, 25 - S7A
* 26 - S8A, 11 - S1B,10 - S2B, 9 - S3B, 8 - S4B, 7 - S5B, 6 - S6B
* 5 - S7B, 4 - S8B, 15 - A2, 16 - A1, 17 - A0, 18 - EN
* 28 - DA, 2 - DB, 1 - VDD, 12 - GND, 27 - VSS
*                    
.SUBCKT ADG407B 19 20 21 22 23 24 25 26 11 10 9 8 7 6 5 4 15 16 17 18 28 2 1 12 27
*
* DEMUX SWITCHES (S1-8A ---> DA) and (S1-8B ---> DB)
*
*     First Section is for control line A0
*          All nodes in this section are in the 30's unless
*          they are I/O nodes
*
E_A0_2    200 12  17 12    1
E_A0_1     30 40 201 40   -1
R_A0_1    200 201         1000
C_A0_X2   201 12          100E-12

V_AX_1     40  12          1.6

SB_A0_8      4 31 201 12  Sdemux
SB_A0_7      5 31 30  12  Sdemux                
SB_A0_6      6 32 201 12  Sdemux
SB_A0_5      7 32 30  12  Sdemux
SB_A0_4      8 33 201 12  Sdemux
SB_A0_3      9 33 30  12  Sdemux
SB_A0_2     10 34 201 12  Sdemux
SB_A0_1     11 34 30  12  Sdemux

SA_A0_8     26 35 201 12  Sdemux
SA_A0_7     25 35 30  12  Sdemux                
SA_A0_6     24 36 201 12  Sdemux
SA_A0_5     23 36 30  12  Sdemux
SA_A0_4     22 37 201 12  Sdemux
SA_A0_3     21 37 30  12  Sdemux
SA_A0_2     20 38 201 12  Sdemux
SA_A0_1     19 38 30  12  Sdemux

CA_A0_X1     17 12          4E-12
CA_A0_D      17 48          4E-12
CB_A0_X1     17 12          4E-12
CB_A0_D      17 47          4E-12

*          Input capacitances

CA_A0_1     19  12         8E-12
CA_A0_2     20  12         8E-12
CA_A0_3     21  12         8E-12
CA_A0_4     22  12         8E-12
CA_A0_5     23  12         8E-12
CA_A0_6     24  12         8E-12
CA_A0_7     25  12         8E-12
CA_A0_8     26  12         8E-12

CB_A0_1    11  12         8E-12
CB_A0_2    10  12         8E-12
CB_A0_3     9  12         8E-12
CB_A0_4     8  12         8E-12
CB_A0_5     7  12         8E-12
CB_A0_6     6  12         8E-12
CB_A0_7     5  12         8E-12
CB_A0_8     4  12         8E-12

C_D_1      28  12         80E-12
C_D_2       2  12         80E-12
*
*       Leakage Current (SX and D ON only) 
*

RA_ON_S1   19 500    12E9
RA_ON_S2   20 500    12E9
RA_ON_S3   21 500    12E9
RA_ON_S4   22 500    12E9
RA_ON_S5   23 500    12E9
RA_ON_S6   24 500    12E9
RA_ON_S7   25 500    12E9
RA_ON_S8   26 500    12E9

RB_ON_S1   11 500    12E9
RB_ON_S2   10 500    12E9
RB_ON_S3    9 500    12E9
RB_ON_S4    8 500    12E9
RB_ON_S5    7 500    12E9
RB_ON_S6    6 500    12E9
RB_ON_S7    5 500    12E9
RB_ON_S8    4 500    12E9

SLEAK_ON_DA 28 500    28 500  SLEAK
ILEAK_ON_DA 28 500    200E-12              

SLEAK_ON_DB 2 500    2 500  SLEAK
ILEAK_ON_DB 2 500    200E-12     
*
*       Leakage Current (SX OFF only)
*
*       Leakage Current (D OFF only)
*

SA_OFF_D     28  58 80 12         Sdemux
RA_OFF_D     58  12                1E12 
GA_OFF_D     28  12 58 12          0.75E-12

SB_OFF_D     2  58 80 12          Sdemux
RB_OFF_D     58  12                1E12 
GB_OFF_D     2  12 58 12          0.75E-12

*
*     Second Section is for control line A1
*

E_A1_2    170 12 16  12    1
E_A1_1     41 40 171 40   -1
R_A1_1    170 171         1000
C_A1_X2   171 12          100E-12

SB_A1_1     31 42 171 12     Sdemux
SB_A1_2     32 42 41  12     Sdemux
SB_A1_3     33 43 171 12    Sdemux
SB_A1_4     34 43 41  12    Sdemux

SA_A1_1     35 44 171 12    Sdemux
SA_A1_2     36 44 41  12    Sdemux
SA_A1_3     37 45 171 12    Sdemux
SA_A1_4     38 45 41  12    Sdemux

CA_A1_X     16 12           4E-12
CA_A1_D     16 48           4E-12
CB_A1_X     16 12           4E-12
CB_A1_D     16 47           4E-12
*
*     Third Section is for control line A2
*

E_A2_2    160 12 15  12    1
E_A2_1     46 40 161 40   -1
R_A2_1    160 161         1000
C_A2_X2   161  12          100E-12

SB_A2_1     42 47 161 12     Sdemux
SB_A2_2     43 47 46  12    Sdemux

SA_A2_3     44 48 161 12    Sdemux
SA_A2_4     45 48 46  12    Sdemux

CA_A2_X     15 12           4E-12
CA_A2_D     15 48           4E-12

CB_A2_X     15 12           4E-12
CB_A2_D     15 47           4E-12

*
*     Main Series Switch combination - A
*
*

VA_1_A     519 500         15
VA_1_B     520 500         -15
RVA_1_A   519 500  1E6
RVA_1_B   520 500 1E6
VA_1_C     521 500         -0.5 ;sets pos main offset
VA_1_D     522  27         2.5  ;sets neg main offset
RA_1_C     48    0         1E13
SA_1_A     525  48 520  83 SNCM
RA_1_A     512 525         24           ;sets neg at max d
SA_1_B     526  48 519  83 SPCM
RA_1_B      83 526         30           ;sets pos at max d
SA_1_C      83 512 711 500 SMAINP
SA_1_D     512 511 500 712 SMAINN
EA_1_E     711 500         VALUE = {(10*V(83,521))/(0.5*V(1,500)+0.005)}
EA_1_F     712 500         VALUE = {(10*V(83,500))/(PWR(V(500,522),1)+0.005)}
SA_1_G     511  48   1  27 SBASE
R_VA_B     521 500 1E6     
R_VA_C     522 500 1E6



*
*     Main Series Switch combination - B
*

VB_1_A     419 500         15
VB_1_B     420 500         -15
RVB_1_A   419 500  1E6
RVB_1_B   420 500 1E6
VB_1_C     421 500         -0.5         ;sets pos main offset
VB_1_D     422  27         2.5          ;sets neg main offset
RB_1_C      47   0         1E13
SB_1_A     425  47 420  73 SNCM
RB_1_A     412 425         24           ;sets neg at max d
SB_1_B     426  47 419  73 SPCM
RB_1_B      73 426         30           ;sets pos at max d
SB_1_C      73 412 611 500 SMAINP
SB_1_D     412 411 500 612 SMAINN
EB_1_E     611 500         VALUE = {(10*V(73,421))/(0.5*V(1,500)+0.005)}
EB_1_F     612 500         VALUE = {(10*V(73,500))/(PWR(V(500,422),1)+0.005)}
SB_1_G     411  47   1  27 SBASE
R_VB_B     421 500 1E6     ;Add dummy resistors so that SPICE has two 
R_VB_C     422 500 1E6             components on these nodes
*
*       Voltage Clamp 
*

DA_1_POS     48  1    DClamp
GA_1_POS     48  1  48  1  -1E-12
DA_2_NEG     27  48   DClamp
GA_2_NEG     27  48 27  48 1E-12

DB_1_POS     47  1    DClamp
GB_1_POS     47  1  47  1  -1E-12
DB_2_NEG     27  47   DClamp
GB_2_NEG     27  47 27  47 1E-12

*     Enable Switch section
*

SB_EN_1     73 2 18  12     Sdemux
SA_EN_1     83  28 18  12     sdemux
CA_EN_1     18  2           4.2E-12
CB_EN_1     18 28           4.2E-12  ; SETS CHARGE INJECTION 

*     Invert Enable Switch section

E_EN0_1     18  81 80 12    -2
V_EN0_1     82  12          2.5
R_EN0_1     82  81         1
R_EN0_2     80  12          1E12

*
*     Power Supply Current Correction
*
I_PS_1      1  12           80E-6
I_PS_2     12  27           0.0001E-6
E_PS_1     99  12  1  12    1
E_PS_2    500  27  1  27    .5
I_E_PS1  99  12  0
*
*       Crosstalk 
*

RAXT_1     19 52           1E13
RAXT_2     20 52           1E13
RAXT_3     21 52           1E13
RAXT_4     22 52           1E13
RAXT_5     23 52           1E13
RAXT_6     24 52           1E13
RAXT_7     25 52           1E13
RAXT_8     26 52           1E13
RBXT_1     11 53           1E13
RBXT_2     10 53           1E13
RBXT_3      9 53           1E13
RBXT_4      8 53           1E13
RBXT_5      7 53           1E13
RBXT_6      6 53           1E13
RBXT_7      5 53           1E13
RBXT_8      4 53           1E13

CAXT_1     19 52           1E-12
CAXT_2     20 52           1E-12
CAXT_3     21 52           1E-12
CAXT_4     22 52           1E-12
CAXT_5     23 52           1E-12
CAXT_6     24 52           1E-12
CAXT_7     25 52           1E-12
CAXT_8     26 52           1E-12

CBXT_1     11 53           1E-12
CBXT_2     10 53           1E-12
CBXT_3      9 53           1E-12
CBXT_4      8 53           1E-12
CBXT_5      7 53           1E-12
CBXT_6      6 53           1E-12
CBXT_7      5 53           1E-12
CBXT_8      4 53           1E-12

*
*       OFF Isolation
*
CAOI_1     19 28           1E-13
CAOI_2     20 28           1E-13
CAOI_3     21 28           1E-13
CAOI_4     22 28           1E-13
CAOI_5     23 28           1E-13
CAOI_6     24 28           1E-13
CAOI_7     25 28           1E-13
CAOI_8     26 28           1E-13
CBOI_9     11  2           1E-13
CBOI_10    10  2           1E-13
CBOI_11     9  2           1E-13
CBOI_12     8  2           1E-13
CBOI_13     7  2           1E-13
CBOI_14     6  2           1E-13
CBOI_15     5  2           1E-13
CBOI_16     4  2           1E-13
RAOI_1     19 1901         1.6E9
CAOI_1A    1901 28         10E-12
RAOI_2     20 1902         1.6E9
CAOI_2A    1902 28         10E-12
RAOI_3     21 1903         1.6E9
CAOI_3A    1903 28         10E-12
RAOI_4     22 1904         1.6E9
CAOI_4A    1904 28         10E-12
RAOI_5     23 1905         1.6E9
CAOI_5A    1905 28         10E-12
RAOI_6     24 1906         1.6E9
CAOI_6A    1906 28         10E-12
RAOI_7     25 1907         1.6E9
CAOI_7A    1907 28         10E-12
RAOI_8     26 1908         1.6E9
CAOI_8A    1908 28         10E-12

RBOI_1     11 1909         1.6E9
CBAOI_1A    1909 2         10E-12
RBOI_2     10 1910         1.6E9
CBOI_2A    1910 2         10E-12
RBOI_3     9 1911         1.6E9
CBOI_3A    1911 2         10E-12
RBOI_4     8 1912         1.6E9
CBOI_4A    1912 2         10E-12
RBOI_5     7 1913         1.6E9
CBOI_5A    1913 2         10E-12
RBOI_6     6 1914         1.6E9
CBOI_6A    1914 2         10E-12
RBOI_7     5 1915         1.6E9
CBOI_7A    1915 2         10E-12
RBOI_8     4 1916         1.6E9
CBOI_8A    1916 2         10E-12
*
* MODELS USED
*
.MODEL SNCM  VSWITCH (RON=30 ROFF=500001 VON=9 VOFF=-44)
.MODEL SPCM  VSWITCH (RON=450000 ROFF=30 VON=41 VOFF=-6.5)
.MODEL SBASE VSWITCH (RON=75 ROFF=3500 VON=28 VOFF=-10)
.MODEL SMAINP VSWITCH (RON=650001 ROFF=60 VON=32 VOFF=0)
.MODEL SMAINN VSWITCH (RON=700001 ROFF=40 VON=28.5 VOFF=0)
.MODEL Sdemux VSWITCH (RON=1 ROFF=1E12 VON=2.0 VOFF=1.4)
.MODEL DClamp D(IS=1E-15 IBV=1E-13)
.MODEL SLEAK VSWITCH (RON=9E8 ROFF=8E8 VON=-15 VOFF=15)
.ENDS ADG407B
