* AD8517/AD8527 SPICE Macro-model
* Typical Values
* 11/99, Ver. 1
* Troy Murphy / ADSC
*
* Copyright 1996 by Analog Devices
*
* Refer to "README.DOC" file for License Statement.  Use of this model
* indicates your acceptance of the terms and provisions in the License
* Statement.
*
* Node Assignments
*			noninverting input
*			|	inverting input
*			|	|	positive supply
*			|	|	|	negative supply
*			|	|	|	|	output
*			|	|	|	|	|
*			|	|	|	|	|
..SUBCKT AD8517	1	2	99	50	45
*
* RAIL-TO-RAIL INPUT STAGE
*
Q1    5  7 3 PIX
Q2    6  2 4 PIX
RC1   5 50 1780
RC2   6 50 1780
RE1   3 10 522
RE2   4 10 522
RCM1 10 99 1.15E+6
CCM1 10 99 3.08E-12
C1    5  6 2.9E-12
D1    3  8 DX
D2    4  9 DX
V1   99  8 DC 0.7
V2   99  9 DC 0.7
I1   99 10 225E-6
Q3   11  7 13 NIX
Q4   12  2 14 NIX
RC3  99 11 1780
RC4  99 12 1780
RE3  13 15 522
RE4  14 15 522
RCM2 15 50 1.15E+6
CCM2 15 50 3.08E-12
C2   11 12 2.9E-12
I2   15 50 225E-6
V3   16 50 DC 0.7
V4   17 50 DC 0.7
D3   16 13 DX
D4   17 14 DX
EOS   7  1 POLY(2) (73,98) (81,98) 1.3E-3 1 1
IOS   1  2 50E-9
*
* PSRR=90dB, ZERO AT 100Hz
*
RPS1 70  0 1E+6
RPS2 71  0 1E+6
CPS1 99 70 1E-5
CPS2 50 71 1E-5
EPSY 98 72 POLY(2) (70,0) (0,71) 0 1 1
RPS3 72 73 15.9E+6
CPS3 72 73 50E-12
RPS4 73 98 480
*
* VOLTAGE NOISE REFERENCE OF 12nV/rt(Hz)
*
VN1 80 98 0
RN1 80 98 16.45E-3
HN  81 98 VN1 12
RN2 81 98 1
*
* INTERNAL VOLTAGE REFERENCE
*
EREF 98  0 POLY(2) (99,0) (50,0) 0 .5 .5
GSY  99 50 POLY(1) (99,50) 56.1E-6 25E-6
EVP  97 98 (99,50) 0.5
EVN  51 98 (50,99) 0.5
*
* GAIN STAGE
*
G1   98 30 POLY(2) (5,6) (11,12) 0 0.8E-3 0.8E-3
R1   30 98 3.47E+5
CF   30 45 80E-12
D5   30 97 DX
D6   51 30 DX
*
* RAIL-TO-RAIL OUTPUT STAGE
*
Q5   45 41 99 POUT
Q6   45 43 50 NOUT
EB1  99 40 POLY(1) (98,30) 0.7308 1
EB2  42 50 POLY(1) (30,98) 0.7308 1
RB1  40 41 500
RB2  42 43 500
D7   46 99 DX
D8   47 43 DX
V5   46 41 0.5
V6   47 50 0.5
*
..MODEL NIX NPN (BF=280,IS=1E-16,VAF=130,KF=2.5E-14)
..MODEL PIX PNP (BF=560,IS=1E-16,VAF=130,KF=2.5E-14)
..MODEL POUT PNP (BF=100,IS=1E-16,VAF=130,RC=20)
..MODEL NOUT NPN (BF=100,IS=1E-16,VAF=130,RC=11)
..MODEL DX D(IS=1E-16,RS=5)
..ENDS AD8517
