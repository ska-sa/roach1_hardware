* AD828 SPICE Model                     Rev. A, 4/93
*                                       ARG / PMI
*
* Copyright 1993 by Analog Devices
*
* Refer to "README.DOC" file for License Statement.  Use of
* this model indicates your acceptance of the terms and pro-
* visions in the License Statement.
*
* Node assignments
*                non-inverting input
*                |  inverting input
*                |  |  positive supply
*                |  |  |  negative supply
*                |  |  |  |  output
*                |  |  |  |  |
.SUBCKT AD828    2  1  99 50 46
*
* INPUT STAGE AND POLE AT 500MHZ
*
I1   4    50   1E-3
CIN  1    2    1.5E-12
CC1  1    0    .5E-12
CC2  2    0    .5E-12
IOS  2    1    25E-9
Q1   5    1    7    QN
Q2   6    3    8    QN
R3   99   5    884
R4   99   6    884
R5   7    4    832
R6   8    4    832
C1   5    6    180E-15
EOS  3    2    POLY(1) (21,98) 500E-6 0.1
*
* GAIN STAGE AND DOMINANT POLE AT 10KHZ
*
EREF 98   0    (39,0) 1
G1   98   9    (5,6) 1.131E-3
R7   9    98   7.958E6
C2   9    98   2E-12
D1   9    10   DX
D2   11   9    DX
V1   99   10   1.8
V2   11   50   1.8
*
* NEGATIVE ZERO AT 150MHZ
*
E1   14   98   (9,39) 1E6
R11  14   15   1
R12  15   98   1E-6
FNZ  14   15   VNZ -1
ENZ  16   98   (14,15) 1
VNZ  17   98   DC 0
CNZ  16   17   1.061E-9
*
* ZERO/POLE AT 60MHZ/75MHZ
*
E2   18   98   (15,39) 1.25
R13  18   19   1
R14  19   98   4
C5   18   19   2.653E-9
*
* COMMON MODE GAIN STAGE WITH ZERO AT 100HZ
*
ECM  20   98   POLY(2) (1,39) (2,39) 0 0.5 0.5
R8   20   21   1E6
R9   21   98   10
C3   20   21   1.592E-9
*
* POLE AT 400MHZ
*
G2   98   40   (19,39) 1E-6
R10  40   98   1E6
C4   40   98   .398E-15
*
* OUTPUT STAGE
*
RS1  99   39   65E3
RS2  39   50   65E3
RO1  99   45   16
RO2  45   50   16
G7   45   99   (99,40) 62.5E-3
G8   50   45   (40,50) 62.5E-3
G9   98   60   (45,40) 62.5E-3
D7   60   61   DX
D8   62   60   DX
V7   61   98   DC 0
V8   98   62   DC 0
FSY  99   50   POLY(2) V7 V8 5.77E-3 1 1
D9   41   45   DX
D10  45   42   DX
V5   40   41   0.4
V6   42   40   0.4
LO   45   46   5E-8
.MODEL QN NPN(BF=150.52)
.MODEL DX D(IS=1E-12)
.ENDS AD828