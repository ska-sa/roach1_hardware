* OP183G SPICE Macro-model              Rev. A, 3/94
*                                       ARG / PMI
*
* This version of the OP183 model simulates the worst-case
* parameters of the 'G' grade.  The worst-case parameters
* used correspond to those in the data sheet.
*
* Copyright 1993 by Analog Devices
*
* Refer to "README.DOC" file for License Statement. Use of
* this model indicates your acceptance of the terms and pro-
* visions in the License Statement.
*
* Node assignments
*                non-inverting input
*                |  inverting input
*                |  |  positive supply
*                |  |  |  negative supply
*                |  |  |  |  output
*                |  |  |  |  |
.SUBCKT OP183G   2  1  99 50 45
*
* INPUT STAGE AND POLE AT 600KHZ
*
I1   99   8    1E-4
Q1   4    1    6    QP
Q2   5    3    7    QP
CIN  1    2    1.5PF
R1   50   4    796
R2   50   5    796
C1   4    5    167E-12
R3   6    8    279
R4   7    8    279
IOS  1    2    25E-9
EOS  3    2    POLY(1) (15,98) 1E-3 1
DC1  2   36    DZ
DC2  1   36    DZ
*
* GAIN STAGE AND DOMINANT POLE AT 100HZ
*
EREF 98   0    POLY(2) (99,0) (50,0) 0 0.5 0.5
G1   98   9    (4,5) 1.257E-3
R5   9    98   79.577E6
C2   9    98   20E-12
D1   9    10   DX
D2   11   9    DX
E1   10   98   POLY(1)  99  98  -1.6185  1.0623
V2   50   11   -0.666
*
* COMMON MODE STAGE WITH ZERO AT 17.7KHZ
*
ECM  14   98   POLY(2) (1,98) (2,98) 0 158 158
R7   14   15   1E6
C4   14   15   9E-12
R8   15   98   1
*
* POLE AT 20MHZ
*
GP2  98   31   (9,98) 1E-6
RP2  31   98   1E6
CP2  31   98   7.96E-15
*
* ZERO AT 1.5MHZ
*
EZ1  32   98   (31,98) 1E6
RZ1  32   33   1E6   
RZ2  33   98   1
CZ1  32   33   106E-15
*
* POLE AT 10MHZ
*
GP10  98   40   (33,98) 1E-6
RP10  40   98   1E6
CP10  40   98   15.9E-15
*
* OUTPUT STAGE
*
RO1  99   45   140
RO2  45   50   140
G7   45   99   (99,40) 7.143E-3
G8   50   45   (40,50) 7.143E-3
G9   98   60   (45,40) 7.143E-3
D7   60   61   DX
D8   62   60   DX
V7   61   98   DC 0
V8   98   62   DC 0
GSY  99   50   (99,50) 5E-6
FSY  99   50   POLY(2) V7 V8 1.375E-3  1  1
D9   40   41   DX
D10  42   40   DX
V5   41   45   1.2
V6   45   42   1.5
*
* MODELS USED
*
.MODEL DX D
.MODEL DZ D(IS=1E-15 BV=7.0)
.MODEL QP PNP(BF=82.333)
.ENDS
